magic
tech sky130B
magscale 1 2
timestamp 1672519886
<< nwell >>
rect 1066 176517 178886 177083
rect 1066 175429 178886 175995
rect 1066 174341 178886 174907
rect 1066 173253 178886 173819
rect 1066 172165 178886 172731
rect 1066 171077 178886 171643
rect 1066 169989 178886 170555
rect 1066 168901 178886 169467
rect 1066 167813 178886 168379
rect 1066 166725 178886 167291
rect 1066 165637 178886 166203
rect 1066 164549 178886 165115
rect 1066 163461 178886 164027
rect 1066 162373 178886 162939
rect 1066 161285 178886 161851
rect 1066 160197 178886 160763
rect 1066 159109 178886 159675
rect 1066 158021 178886 158587
rect 1066 156933 178886 157499
rect 1066 155845 178886 156411
rect 1066 154757 178886 155323
rect 1066 153669 178886 154235
rect 1066 152581 178886 153147
rect 1066 151493 178886 152059
rect 1066 150405 178886 150971
rect 1066 149317 178886 149883
rect 1066 148229 178886 148795
rect 1066 147141 178886 147707
rect 1066 146053 178886 146619
rect 1066 144965 178886 145531
rect 1066 143877 178886 144443
rect 1066 142789 178886 143355
rect 1066 141701 178886 142267
rect 1066 140613 178886 141179
rect 1066 139525 178886 140091
rect 1066 138437 178886 139003
rect 1066 137349 178886 137915
rect 1066 136261 178886 136827
rect 1066 135173 178886 135739
rect 1066 134085 178886 134651
rect 1066 132997 178886 133563
rect 1066 131909 178886 132475
rect 1066 130821 178886 131387
rect 1066 129733 178886 130299
rect 1066 128645 178886 129211
rect 1066 127557 178886 128123
rect 1066 126469 178886 127035
rect 1066 125381 178886 125947
rect 1066 124293 178886 124859
rect 1066 123205 178886 123771
rect 1066 122117 178886 122683
rect 1066 121029 178886 121595
rect 1066 119941 178886 120507
rect 1066 118853 178886 119419
rect 1066 117765 178886 118331
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 177361
<< obsm1 >>
rect 1104 2128 178848 178220
<< metal2 >>
rect 2594 179200 2650 180000
rect 4986 179200 5042 180000
rect 7378 179200 7434 180000
rect 9770 179200 9826 180000
rect 12162 179200 12218 180000
rect 14554 179200 14610 180000
rect 16946 179200 17002 180000
rect 19338 179200 19394 180000
rect 21730 179200 21786 180000
rect 24122 179200 24178 180000
rect 26514 179200 26570 180000
rect 28906 179200 28962 180000
rect 31298 179200 31354 180000
rect 33690 179200 33746 180000
rect 36082 179200 36138 180000
rect 38474 179200 38530 180000
rect 40866 179200 40922 180000
rect 43258 179200 43314 180000
rect 45650 179200 45706 180000
rect 48042 179200 48098 180000
rect 50434 179200 50490 180000
rect 52826 179200 52882 180000
rect 55218 179200 55274 180000
rect 57610 179200 57666 180000
rect 60002 179200 60058 180000
rect 62394 179200 62450 180000
rect 64786 179200 64842 180000
rect 67178 179200 67234 180000
rect 69570 179200 69626 180000
rect 71962 179200 72018 180000
rect 74354 179200 74410 180000
rect 76746 179200 76802 180000
rect 79138 179200 79194 180000
rect 81530 179200 81586 180000
rect 83922 179200 83978 180000
rect 86314 179200 86370 180000
rect 88706 179200 88762 180000
rect 91098 179200 91154 180000
rect 93490 179200 93546 180000
rect 95882 179200 95938 180000
rect 98274 179200 98330 180000
rect 100666 179200 100722 180000
rect 103058 179200 103114 180000
rect 105450 179200 105506 180000
rect 107842 179200 107898 180000
rect 110234 179200 110290 180000
rect 112626 179200 112682 180000
rect 115018 179200 115074 180000
rect 117410 179200 117466 180000
rect 119802 179200 119858 180000
rect 122194 179200 122250 180000
rect 124586 179200 124642 180000
rect 126978 179200 127034 180000
rect 129370 179200 129426 180000
rect 131762 179200 131818 180000
rect 134154 179200 134210 180000
rect 136546 179200 136602 180000
rect 138938 179200 138994 180000
rect 141330 179200 141386 180000
rect 143722 179200 143778 180000
rect 146114 179200 146170 180000
rect 148506 179200 148562 180000
rect 150898 179200 150954 180000
rect 153290 179200 153346 180000
rect 155682 179200 155738 180000
rect 158074 179200 158130 180000
rect 160466 179200 160522 180000
rect 162858 179200 162914 180000
rect 165250 179200 165306 180000
rect 167642 179200 167698 180000
rect 170034 179200 170090 180000
rect 172426 179200 172482 180000
rect 174818 179200 174874 180000
rect 177210 179200 177266 180000
rect 44914 0 44970 800
rect 134890 0 134946 800
<< obsm2 >>
rect 2706 179144 4930 179330
rect 5098 179144 7322 179330
rect 7490 179144 9714 179330
rect 9882 179144 12106 179330
rect 12274 179144 14498 179330
rect 14666 179144 16890 179330
rect 17058 179144 19282 179330
rect 19450 179144 21674 179330
rect 21842 179144 24066 179330
rect 24234 179144 26458 179330
rect 26626 179144 28850 179330
rect 29018 179144 31242 179330
rect 31410 179144 33634 179330
rect 33802 179144 36026 179330
rect 36194 179144 38418 179330
rect 38586 179144 40810 179330
rect 40978 179144 43202 179330
rect 43370 179144 45594 179330
rect 45762 179144 47986 179330
rect 48154 179144 50378 179330
rect 50546 179144 52770 179330
rect 52938 179144 55162 179330
rect 55330 179144 57554 179330
rect 57722 179144 59946 179330
rect 60114 179144 62338 179330
rect 62506 179144 64730 179330
rect 64898 179144 67122 179330
rect 67290 179144 69514 179330
rect 69682 179144 71906 179330
rect 72074 179144 74298 179330
rect 74466 179144 76690 179330
rect 76858 179144 79082 179330
rect 79250 179144 81474 179330
rect 81642 179144 83866 179330
rect 84034 179144 86258 179330
rect 86426 179144 88650 179330
rect 88818 179144 91042 179330
rect 91210 179144 93434 179330
rect 93602 179144 95826 179330
rect 95994 179144 98218 179330
rect 98386 179144 100610 179330
rect 100778 179144 103002 179330
rect 103170 179144 105394 179330
rect 105562 179144 107786 179330
rect 107954 179144 110178 179330
rect 110346 179144 112570 179330
rect 112738 179144 114962 179330
rect 115130 179144 117354 179330
rect 117522 179144 119746 179330
rect 119914 179144 122138 179330
rect 122306 179144 124530 179330
rect 124698 179144 126922 179330
rect 127090 179144 129314 179330
rect 129482 179144 131706 179330
rect 131874 179144 134098 179330
rect 134266 179144 136490 179330
rect 136658 179144 138882 179330
rect 139050 179144 141274 179330
rect 141442 179144 143666 179330
rect 143834 179144 146058 179330
rect 146226 179144 148450 179330
rect 148618 179144 150842 179330
rect 151010 179144 153234 179330
rect 153402 179144 155626 179330
rect 155794 179144 158018 179330
rect 158186 179144 160410 179330
rect 160578 179144 162802 179330
rect 162970 179144 165194 179330
rect 165362 179144 167586 179330
rect 167754 179144 169978 179330
rect 170146 179144 172370 179330
rect 172538 179144 174762 179330
rect 174930 179144 177154 179330
rect 177322 179144 177540 179330
rect 2596 856 177540 179144
rect 2596 800 44858 856
rect 45026 800 134834 856
rect 135002 800 177540 856
<< obsm3 >>
rect 4210 2143 173486 177853
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
<< obsm4 >>
rect 45875 3435 50208 176901
rect 50688 3435 65568 176901
rect 66048 3435 80928 176901
rect 81408 3435 96288 176901
rect 96768 3435 111648 176901
rect 112128 3435 127008 176901
rect 127488 3435 129477 176901
<< labels >>
rlabel metal2 s 167642 179200 167698 180000 6 Dataw_en
port 1 nsew signal output
rlabel metal2 s 174818 179200 174874 180000 6 Serial_input
port 2 nsew signal input
rlabel metal2 s 177210 179200 177266 180000 6 Serial_output
port 3 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 clk
port 4 nsew signal input
rlabel metal2 s 71962 179200 72018 180000 6 data_mem_addr[0]
port 5 nsew signal output
rlabel metal2 s 74354 179200 74410 180000 6 data_mem_addr[1]
port 6 nsew signal output
rlabel metal2 s 76746 179200 76802 180000 6 data_mem_addr[2]
port 7 nsew signal output
rlabel metal2 s 79138 179200 79194 180000 6 data_mem_addr[3]
port 8 nsew signal output
rlabel metal2 s 81530 179200 81586 180000 6 data_mem_addr[4]
port 9 nsew signal output
rlabel metal2 s 83922 179200 83978 180000 6 data_mem_addr[5]
port 10 nsew signal output
rlabel metal2 s 86314 179200 86370 180000 6 data_mem_addr[6]
port 11 nsew signal output
rlabel metal2 s 88706 179200 88762 180000 6 data_mem_addr[7]
port 12 nsew signal output
rlabel metal2 s 172426 179200 172482 180000 6 hlt
port 13 nsew signal output
rlabel metal2 s 2594 179200 2650 180000 6 instr[0]
port 14 nsew signal input
rlabel metal2 s 50434 179200 50490 180000 6 instr[10]
port 15 nsew signal input
rlabel metal2 s 55218 179200 55274 180000 6 instr[11]
port 16 nsew signal input
rlabel metal2 s 60002 179200 60058 180000 6 instr[12]
port 17 nsew signal input
rlabel metal2 s 64786 179200 64842 180000 6 instr[13]
port 18 nsew signal input
rlabel metal2 s 67178 179200 67234 180000 6 instr[14]
port 19 nsew signal input
rlabel metal2 s 69570 179200 69626 180000 6 instr[15]
port 20 nsew signal input
rlabel metal2 s 7378 179200 7434 180000 6 instr[1]
port 21 nsew signal input
rlabel metal2 s 12162 179200 12218 180000 6 instr[2]
port 22 nsew signal input
rlabel metal2 s 16946 179200 17002 180000 6 instr[3]
port 23 nsew signal input
rlabel metal2 s 21730 179200 21786 180000 6 instr[4]
port 24 nsew signal input
rlabel metal2 s 26514 179200 26570 180000 6 instr[5]
port 25 nsew signal input
rlabel metal2 s 31298 179200 31354 180000 6 instr[6]
port 26 nsew signal input
rlabel metal2 s 36082 179200 36138 180000 6 instr[7]
port 27 nsew signal input
rlabel metal2 s 40866 179200 40922 180000 6 instr[8]
port 28 nsew signal input
rlabel metal2 s 45650 179200 45706 180000 6 instr[9]
port 29 nsew signal input
rlabel metal2 s 4986 179200 5042 180000 6 instr_mem_addr[0]
port 30 nsew signal output
rlabel metal2 s 52826 179200 52882 180000 6 instr_mem_addr[10]
port 31 nsew signal output
rlabel metal2 s 57610 179200 57666 180000 6 instr_mem_addr[11]
port 32 nsew signal output
rlabel metal2 s 62394 179200 62450 180000 6 instr_mem_addr[12]
port 33 nsew signal output
rlabel metal2 s 9770 179200 9826 180000 6 instr_mem_addr[1]
port 34 nsew signal output
rlabel metal2 s 14554 179200 14610 180000 6 instr_mem_addr[2]
port 35 nsew signal output
rlabel metal2 s 19338 179200 19394 180000 6 instr_mem_addr[3]
port 36 nsew signal output
rlabel metal2 s 24122 179200 24178 180000 6 instr_mem_addr[4]
port 37 nsew signal output
rlabel metal2 s 28906 179200 28962 180000 6 instr_mem_addr[5]
port 38 nsew signal output
rlabel metal2 s 33690 179200 33746 180000 6 instr_mem_addr[6]
port 39 nsew signal output
rlabel metal2 s 38474 179200 38530 180000 6 instr_mem_addr[7]
port 40 nsew signal output
rlabel metal2 s 43258 179200 43314 180000 6 instr_mem_addr[8]
port 41 nsew signal output
rlabel metal2 s 48042 179200 48098 180000 6 instr_mem_addr[9]
port 42 nsew signal output
rlabel metal2 s 91098 179200 91154 180000 6 read_data[0]
port 43 nsew signal input
rlabel metal2 s 115018 179200 115074 180000 6 read_data[10]
port 44 nsew signal input
rlabel metal2 s 117410 179200 117466 180000 6 read_data[11]
port 45 nsew signal input
rlabel metal2 s 119802 179200 119858 180000 6 read_data[12]
port 46 nsew signal input
rlabel metal2 s 122194 179200 122250 180000 6 read_data[13]
port 47 nsew signal input
rlabel metal2 s 124586 179200 124642 180000 6 read_data[14]
port 48 nsew signal input
rlabel metal2 s 126978 179200 127034 180000 6 read_data[15]
port 49 nsew signal input
rlabel metal2 s 93490 179200 93546 180000 6 read_data[1]
port 50 nsew signal input
rlabel metal2 s 95882 179200 95938 180000 6 read_data[2]
port 51 nsew signal input
rlabel metal2 s 98274 179200 98330 180000 6 read_data[3]
port 52 nsew signal input
rlabel metal2 s 100666 179200 100722 180000 6 read_data[4]
port 53 nsew signal input
rlabel metal2 s 103058 179200 103114 180000 6 read_data[5]
port 54 nsew signal input
rlabel metal2 s 105450 179200 105506 180000 6 read_data[6]
port 55 nsew signal input
rlabel metal2 s 107842 179200 107898 180000 6 read_data[7]
port 56 nsew signal input
rlabel metal2 s 110234 179200 110290 180000 6 read_data[8]
port 57 nsew signal input
rlabel metal2 s 112626 179200 112682 180000 6 read_data[9]
port 58 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 reset
port 59 nsew signal input
rlabel metal2 s 170034 179200 170090 180000 6 start
port 60 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 62 nsew ground bidirectional
rlabel metal2 s 129370 179200 129426 180000 6 write_data[0]
port 63 nsew signal output
rlabel metal2 s 153290 179200 153346 180000 6 write_data[10]
port 64 nsew signal output
rlabel metal2 s 155682 179200 155738 180000 6 write_data[11]
port 65 nsew signal output
rlabel metal2 s 158074 179200 158130 180000 6 write_data[12]
port 66 nsew signal output
rlabel metal2 s 160466 179200 160522 180000 6 write_data[13]
port 67 nsew signal output
rlabel metal2 s 162858 179200 162914 180000 6 write_data[14]
port 68 nsew signal output
rlabel metal2 s 165250 179200 165306 180000 6 write_data[15]
port 69 nsew signal output
rlabel metal2 s 131762 179200 131818 180000 6 write_data[1]
port 70 nsew signal output
rlabel metal2 s 134154 179200 134210 180000 6 write_data[2]
port 71 nsew signal output
rlabel metal2 s 136546 179200 136602 180000 6 write_data[3]
port 72 nsew signal output
rlabel metal2 s 138938 179200 138994 180000 6 write_data[4]
port 73 nsew signal output
rlabel metal2 s 141330 179200 141386 180000 6 write_data[5]
port 74 nsew signal output
rlabel metal2 s 143722 179200 143778 180000 6 write_data[6]
port 75 nsew signal output
rlabel metal2 s 146114 179200 146170 180000 6 write_data[7]
port 76 nsew signal output
rlabel metal2 s 148506 179200 148562 180000 6 write_data[8]
port 77 nsew signal output
rlabel metal2 s 150898 179200 150954 180000 6 write_data[9]
port 78 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 24911872
string GDS_FILE /home/radhe/mpw8/caravel_user_project/openlane/processor/runs/23_01_01_02_06/results/signoff/processor.magic.gds
string GDS_START 617782
<< end >>

