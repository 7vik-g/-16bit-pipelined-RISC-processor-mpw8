magic
tech sky130B
magscale 1 2
timestamp 1672520698
<< nwell >>
rect 1066 197189 198850 197510
rect 1066 196101 198850 196667
rect 1066 195013 198850 195579
rect 1066 193925 198850 194491
rect 1066 192837 198850 193403
rect 1066 191749 198850 192315
rect 1066 190661 198850 191227
rect 1066 189573 198850 190139
rect 1066 188485 198850 189051
rect 1066 187397 198850 187963
rect 1066 186309 198850 186875
rect 1066 185221 198850 185787
rect 1066 184133 198850 184699
rect 1066 183045 198850 183611
rect 1066 181957 198850 182523
rect 1066 180869 198850 181435
rect 1066 179781 198850 180347
rect 1066 178693 198850 179259
rect 1066 177605 198850 178171
rect 1066 176517 198850 177083
rect 1066 175429 198850 175995
rect 1066 174341 198850 174907
rect 1066 173253 198850 173819
rect 1066 172165 198850 172731
rect 1066 171077 198850 171643
rect 1066 169989 198850 170555
rect 1066 168901 198850 169467
rect 1066 167813 198850 168379
rect 1066 166725 198850 167291
rect 1066 165637 198850 166203
rect 1066 164549 198850 165115
rect 1066 163461 198850 164027
rect 1066 162373 198850 162939
rect 1066 161285 198850 161851
rect 1066 160197 198850 160763
rect 1066 159109 198850 159675
rect 1066 158021 198850 158587
rect 1066 156933 198850 157499
rect 1066 155845 198850 156411
rect 1066 154757 198850 155323
rect 1066 153669 198850 154235
rect 1066 152581 198850 153147
rect 1066 151493 198850 152059
rect 1066 150405 198850 150971
rect 1066 149317 198850 149883
rect 1066 148229 198850 148795
rect 1066 147141 198850 147707
rect 1066 146053 198850 146619
rect 1066 144965 198850 145531
rect 1066 143877 198850 144443
rect 1066 142789 198850 143355
rect 1066 141701 198850 142267
rect 1066 140613 198850 141179
rect 1066 139525 198850 140091
rect 1066 138437 198850 139003
rect 1066 137349 198850 137915
rect 1066 136261 198850 136827
rect 1066 135173 198850 135739
rect 1066 134085 198850 134651
rect 1066 132997 198850 133563
rect 1066 131909 198850 132475
rect 1066 130821 198850 131387
rect 1066 129733 198850 130299
rect 1066 128645 198850 129211
rect 1066 127557 198850 128123
rect 1066 126469 198850 127035
rect 1066 125381 198850 125947
rect 1066 124293 198850 124859
rect 1066 123205 198850 123771
rect 1066 122117 198850 122683
rect 1066 121029 198850 121595
rect 1066 119941 198850 120507
rect 1066 118853 198850 119419
rect 1066 117765 198850 118331
rect 1066 116677 198850 117243
rect 1066 115589 198850 116155
rect 1066 114501 198850 115067
rect 1066 113413 198850 113979
rect 1066 112325 198850 112891
rect 1066 111237 198850 111803
rect 1066 110149 198850 110715
rect 1066 109061 198850 109627
rect 1066 107973 198850 108539
rect 1066 106885 198850 107451
rect 1066 105797 198850 106363
rect 1066 104709 198850 105275
rect 1066 103621 198850 104187
rect 1066 102533 198850 103099
rect 1066 101445 198850 102011
rect 1066 100357 198850 100923
rect 1066 99269 198850 99835
rect 1066 98181 198850 98747
rect 1066 97093 198850 97659
rect 1066 96005 198850 96571
rect 1066 94917 198850 95483
rect 1066 93829 198850 94395
rect 1066 92741 198850 93307
rect 1066 91653 198850 92219
rect 1066 90565 198850 91131
rect 1066 89477 198850 90043
rect 1066 88389 198850 88955
rect 1066 87301 198850 87867
rect 1066 86213 198850 86779
rect 1066 85125 198850 85691
rect 1066 84037 198850 84603
rect 1066 82949 198850 83515
rect 1066 81861 198850 82427
rect 1066 80773 198850 81339
rect 1066 79685 198850 80251
rect 1066 78597 198850 79163
rect 1066 77509 198850 78075
rect 1066 76421 198850 76987
rect 1066 75333 198850 75899
rect 1066 74245 198850 74811
rect 1066 73157 198850 73723
rect 1066 72069 198850 72635
rect 1066 70981 198850 71547
rect 1066 69893 198850 70459
rect 1066 68805 198850 69371
rect 1066 67717 198850 68283
rect 1066 66629 198850 67195
rect 1066 65541 198850 66107
rect 1066 64453 198850 65019
rect 1066 63365 198850 63931
rect 1066 62277 198850 62843
rect 1066 61189 198850 61755
rect 1066 60101 198850 60667
rect 1066 59013 198850 59579
rect 1066 57925 198850 58491
rect 1066 56837 198850 57403
rect 1066 55749 198850 56315
rect 1066 54661 198850 55227
rect 1066 53573 198850 54139
rect 1066 52485 198850 53051
rect 1066 51397 198850 51963
rect 1066 50309 198850 50875
rect 1066 49221 198850 49787
rect 1066 48133 198850 48699
rect 1066 47045 198850 47611
rect 1066 45957 198850 46523
rect 1066 44869 198850 45435
rect 1066 43781 198850 44347
rect 1066 42693 198850 43259
rect 1066 41605 198850 42171
rect 1066 40517 198850 41083
rect 1066 39429 198850 39995
rect 1066 38341 198850 38907
rect 1066 37253 198850 37819
rect 1066 36165 198850 36731
rect 1066 35077 198850 35643
rect 1066 33989 198850 34555
rect 1066 32901 198850 33467
rect 1066 31813 198850 32379
rect 1066 30725 198850 31291
rect 1066 29637 198850 30203
rect 1066 28549 198850 29115
rect 1066 27461 198850 28027
rect 1066 26373 198850 26939
rect 1066 25285 198850 25851
rect 1066 24197 198850 24763
rect 1066 23109 198850 23675
rect 1066 22021 198850 22587
rect 1066 20933 198850 21499
rect 1066 19845 198850 20411
rect 1066 18757 198850 19323
rect 1066 17669 198850 18235
rect 1066 16581 198850 17147
rect 1066 15493 198850 16059
rect 1066 14405 198850 14971
rect 1066 13317 198850 13883
rect 1066 12229 198850 12795
rect 1066 11141 198850 11707
rect 1066 10053 198850 10619
rect 1066 8965 198850 9531
rect 1066 7877 198850 8443
rect 1066 6789 198850 7355
rect 1066 5701 198850 6267
rect 1066 4613 198850 5179
rect 1066 3525 198850 4091
rect 1066 2437 198850 3003
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 1104 1980 198812 199436
<< metal2 >>
rect 3698 199200 3754 200000
rect 4066 199200 4122 200000
rect 4434 199200 4490 200000
rect 4802 199200 4858 200000
rect 5170 199200 5226 200000
rect 5538 199200 5594 200000
rect 5906 199200 5962 200000
rect 6274 199200 6330 200000
rect 6642 199200 6698 200000
rect 7010 199200 7066 200000
rect 7378 199200 7434 200000
rect 7746 199200 7802 200000
rect 8114 199200 8170 200000
rect 8482 199200 8538 200000
rect 8850 199200 8906 200000
rect 9218 199200 9274 200000
rect 9586 199200 9642 200000
rect 9954 199200 10010 200000
rect 10322 199200 10378 200000
rect 10690 199200 10746 200000
rect 11058 199200 11114 200000
rect 11426 199200 11482 200000
rect 11794 199200 11850 200000
rect 12162 199200 12218 200000
rect 12530 199200 12586 200000
rect 12898 199200 12954 200000
rect 13266 199200 13322 200000
rect 13634 199200 13690 200000
rect 14002 199200 14058 200000
rect 14370 199200 14426 200000
rect 14738 199200 14794 200000
rect 15106 199200 15162 200000
rect 15474 199200 15530 200000
rect 15842 199200 15898 200000
rect 16210 199200 16266 200000
rect 16578 199200 16634 200000
rect 16946 199200 17002 200000
rect 17314 199200 17370 200000
rect 17682 199200 17738 200000
rect 18050 199200 18106 200000
rect 18418 199200 18474 200000
rect 18786 199200 18842 200000
rect 19154 199200 19210 200000
rect 19522 199200 19578 200000
rect 19890 199200 19946 200000
rect 20258 199200 20314 200000
rect 20626 199200 20682 200000
rect 20994 199200 21050 200000
rect 21362 199200 21418 200000
rect 21730 199200 21786 200000
rect 22098 199200 22154 200000
rect 22466 199200 22522 200000
rect 22834 199200 22890 200000
rect 23202 199200 23258 200000
rect 23570 199200 23626 200000
rect 23938 199200 23994 200000
rect 24306 199200 24362 200000
rect 24674 199200 24730 200000
rect 25042 199200 25098 200000
rect 25410 199200 25466 200000
rect 25778 199200 25834 200000
rect 26146 199200 26202 200000
rect 26514 199200 26570 200000
rect 26882 199200 26938 200000
rect 27250 199200 27306 200000
rect 27618 199200 27674 200000
rect 27986 199200 28042 200000
rect 28354 199200 28410 200000
rect 28722 199200 28778 200000
rect 29090 199200 29146 200000
rect 29458 199200 29514 200000
rect 29826 199200 29882 200000
rect 30194 199200 30250 200000
rect 30562 199200 30618 200000
rect 30930 199200 30986 200000
rect 31298 199200 31354 200000
rect 31666 199200 31722 200000
rect 32034 199200 32090 200000
rect 32402 199200 32458 200000
rect 32770 199200 32826 200000
rect 33138 199200 33194 200000
rect 33506 199200 33562 200000
rect 33874 199200 33930 200000
rect 34242 199200 34298 200000
rect 34610 199200 34666 200000
rect 34978 199200 35034 200000
rect 35346 199200 35402 200000
rect 35714 199200 35770 200000
rect 36082 199200 36138 200000
rect 36450 199200 36506 200000
rect 36818 199200 36874 200000
rect 37186 199200 37242 200000
rect 37554 199200 37610 200000
rect 37922 199200 37978 200000
rect 38290 199200 38346 200000
rect 38658 199200 38714 200000
rect 39026 199200 39082 200000
rect 39394 199200 39450 200000
rect 39762 199200 39818 200000
rect 40130 199200 40186 200000
rect 40498 199200 40554 200000
rect 40866 199200 40922 200000
rect 41234 199200 41290 200000
rect 41602 199200 41658 200000
rect 41970 199200 42026 200000
rect 42338 199200 42394 200000
rect 42706 199200 42762 200000
rect 43074 199200 43130 200000
rect 43442 199200 43498 200000
rect 43810 199200 43866 200000
rect 44178 199200 44234 200000
rect 44546 199200 44602 200000
rect 44914 199200 44970 200000
rect 45282 199200 45338 200000
rect 45650 199200 45706 200000
rect 46018 199200 46074 200000
rect 46386 199200 46442 200000
rect 46754 199200 46810 200000
rect 47122 199200 47178 200000
rect 47490 199200 47546 200000
rect 47858 199200 47914 200000
rect 48226 199200 48282 200000
rect 48594 199200 48650 200000
rect 48962 199200 49018 200000
rect 49330 199200 49386 200000
rect 49698 199200 49754 200000
rect 50066 199200 50122 200000
rect 50434 199200 50490 200000
rect 50802 199200 50858 200000
rect 51170 199200 51226 200000
rect 51538 199200 51594 200000
rect 51906 199200 51962 200000
rect 52274 199200 52330 200000
rect 52642 199200 52698 200000
rect 53010 199200 53066 200000
rect 53378 199200 53434 200000
rect 53746 199200 53802 200000
rect 54114 199200 54170 200000
rect 54482 199200 54538 200000
rect 54850 199200 54906 200000
rect 55218 199200 55274 200000
rect 55586 199200 55642 200000
rect 55954 199200 56010 200000
rect 56322 199200 56378 200000
rect 56690 199200 56746 200000
rect 57058 199200 57114 200000
rect 57426 199200 57482 200000
rect 57794 199200 57850 200000
rect 58162 199200 58218 200000
rect 58530 199200 58586 200000
rect 58898 199200 58954 200000
rect 59266 199200 59322 200000
rect 59634 199200 59690 200000
rect 60002 199200 60058 200000
rect 60370 199200 60426 200000
rect 60738 199200 60794 200000
rect 61106 199200 61162 200000
rect 61474 199200 61530 200000
rect 61842 199200 61898 200000
rect 62210 199200 62266 200000
rect 62578 199200 62634 200000
rect 62946 199200 63002 200000
rect 63314 199200 63370 200000
rect 63682 199200 63738 200000
rect 64050 199200 64106 200000
rect 64418 199200 64474 200000
rect 64786 199200 64842 200000
rect 65154 199200 65210 200000
rect 65522 199200 65578 200000
rect 65890 199200 65946 200000
rect 66258 199200 66314 200000
rect 66626 199200 66682 200000
rect 66994 199200 67050 200000
rect 67362 199200 67418 200000
rect 67730 199200 67786 200000
rect 68098 199200 68154 200000
rect 68466 199200 68522 200000
rect 68834 199200 68890 200000
rect 69202 199200 69258 200000
rect 69570 199200 69626 200000
rect 69938 199200 69994 200000
rect 70306 199200 70362 200000
rect 70674 199200 70730 200000
rect 71042 199200 71098 200000
rect 71410 199200 71466 200000
rect 71778 199200 71834 200000
rect 72146 199200 72202 200000
rect 72514 199200 72570 200000
rect 72882 199200 72938 200000
rect 73250 199200 73306 200000
rect 73618 199200 73674 200000
rect 73986 199200 74042 200000
rect 74354 199200 74410 200000
rect 74722 199200 74778 200000
rect 75090 199200 75146 200000
rect 75458 199200 75514 200000
rect 75826 199200 75882 200000
rect 76194 199200 76250 200000
rect 76562 199200 76618 200000
rect 76930 199200 76986 200000
rect 77298 199200 77354 200000
rect 77666 199200 77722 200000
rect 78034 199200 78090 200000
rect 78402 199200 78458 200000
rect 78770 199200 78826 200000
rect 79138 199200 79194 200000
rect 79506 199200 79562 200000
rect 79874 199200 79930 200000
rect 80242 199200 80298 200000
rect 80610 199200 80666 200000
rect 80978 199200 81034 200000
rect 81346 199200 81402 200000
rect 81714 199200 81770 200000
rect 82082 199200 82138 200000
rect 82450 199200 82506 200000
rect 82818 199200 82874 200000
rect 83186 199200 83242 200000
rect 83554 199200 83610 200000
rect 83922 199200 83978 200000
rect 84290 199200 84346 200000
rect 84658 199200 84714 200000
rect 85026 199200 85082 200000
rect 85394 199200 85450 200000
rect 85762 199200 85818 200000
rect 86130 199200 86186 200000
rect 86498 199200 86554 200000
rect 86866 199200 86922 200000
rect 87234 199200 87290 200000
rect 87602 199200 87658 200000
rect 87970 199200 88026 200000
rect 88338 199200 88394 200000
rect 88706 199200 88762 200000
rect 89074 199200 89130 200000
rect 89442 199200 89498 200000
rect 89810 199200 89866 200000
rect 90178 199200 90234 200000
rect 90546 199200 90602 200000
rect 90914 199200 90970 200000
rect 91282 199200 91338 200000
rect 91650 199200 91706 200000
rect 92018 199200 92074 200000
rect 92386 199200 92442 200000
rect 92754 199200 92810 200000
rect 93122 199200 93178 200000
rect 93490 199200 93546 200000
rect 93858 199200 93914 200000
rect 94226 199200 94282 200000
rect 94594 199200 94650 200000
rect 94962 199200 95018 200000
rect 95330 199200 95386 200000
rect 95698 199200 95754 200000
rect 96066 199200 96122 200000
rect 96434 199200 96490 200000
rect 96802 199200 96858 200000
rect 97170 199200 97226 200000
rect 97538 199200 97594 200000
rect 97906 199200 97962 200000
rect 98274 199200 98330 200000
rect 98642 199200 98698 200000
rect 99010 199200 99066 200000
rect 99378 199200 99434 200000
rect 99746 199200 99802 200000
rect 100114 199200 100170 200000
rect 100482 199200 100538 200000
rect 100850 199200 100906 200000
rect 101218 199200 101274 200000
rect 101586 199200 101642 200000
rect 101954 199200 102010 200000
rect 102322 199200 102378 200000
rect 102690 199200 102746 200000
rect 103058 199200 103114 200000
rect 103426 199200 103482 200000
rect 103794 199200 103850 200000
rect 104162 199200 104218 200000
rect 104530 199200 104586 200000
rect 104898 199200 104954 200000
rect 105266 199200 105322 200000
rect 105634 199200 105690 200000
rect 106002 199200 106058 200000
rect 106370 199200 106426 200000
rect 106738 199200 106794 200000
rect 107106 199200 107162 200000
rect 107474 199200 107530 200000
rect 107842 199200 107898 200000
rect 108210 199200 108266 200000
rect 108578 199200 108634 200000
rect 108946 199200 109002 200000
rect 109314 199200 109370 200000
rect 109682 199200 109738 200000
rect 110050 199200 110106 200000
rect 110418 199200 110474 200000
rect 110786 199200 110842 200000
rect 111154 199200 111210 200000
rect 111522 199200 111578 200000
rect 111890 199200 111946 200000
rect 112258 199200 112314 200000
rect 112626 199200 112682 200000
rect 112994 199200 113050 200000
rect 113362 199200 113418 200000
rect 113730 199200 113786 200000
rect 114098 199200 114154 200000
rect 114466 199200 114522 200000
rect 114834 199200 114890 200000
rect 115202 199200 115258 200000
rect 115570 199200 115626 200000
rect 115938 199200 115994 200000
rect 116306 199200 116362 200000
rect 116674 199200 116730 200000
rect 117042 199200 117098 200000
rect 117410 199200 117466 200000
rect 117778 199200 117834 200000
rect 118146 199200 118202 200000
rect 118514 199200 118570 200000
rect 118882 199200 118938 200000
rect 119250 199200 119306 200000
rect 119618 199200 119674 200000
rect 119986 199200 120042 200000
rect 120354 199200 120410 200000
rect 120722 199200 120778 200000
rect 121090 199200 121146 200000
rect 121458 199200 121514 200000
rect 121826 199200 121882 200000
rect 122194 199200 122250 200000
rect 122562 199200 122618 200000
rect 122930 199200 122986 200000
rect 123298 199200 123354 200000
rect 123666 199200 123722 200000
rect 124034 199200 124090 200000
rect 124402 199200 124458 200000
rect 124770 199200 124826 200000
rect 125138 199200 125194 200000
rect 125506 199200 125562 200000
rect 125874 199200 125930 200000
rect 126242 199200 126298 200000
rect 126610 199200 126666 200000
rect 126978 199200 127034 200000
rect 127346 199200 127402 200000
rect 127714 199200 127770 200000
rect 128082 199200 128138 200000
rect 128450 199200 128506 200000
rect 128818 199200 128874 200000
rect 129186 199200 129242 200000
rect 129554 199200 129610 200000
rect 129922 199200 129978 200000
rect 130290 199200 130346 200000
rect 130658 199200 130714 200000
rect 131026 199200 131082 200000
rect 131394 199200 131450 200000
rect 131762 199200 131818 200000
rect 132130 199200 132186 200000
rect 132498 199200 132554 200000
rect 132866 199200 132922 200000
rect 133234 199200 133290 200000
rect 133602 199200 133658 200000
rect 133970 199200 134026 200000
rect 134338 199200 134394 200000
rect 134706 199200 134762 200000
rect 135074 199200 135130 200000
rect 135442 199200 135498 200000
rect 135810 199200 135866 200000
rect 136178 199200 136234 200000
rect 136546 199200 136602 200000
rect 136914 199200 136970 200000
rect 137282 199200 137338 200000
rect 137650 199200 137706 200000
rect 138018 199200 138074 200000
rect 138386 199200 138442 200000
rect 138754 199200 138810 200000
rect 139122 199200 139178 200000
rect 139490 199200 139546 200000
rect 139858 199200 139914 200000
rect 140226 199200 140282 200000
rect 140594 199200 140650 200000
rect 140962 199200 141018 200000
rect 141330 199200 141386 200000
rect 141698 199200 141754 200000
rect 142066 199200 142122 200000
rect 142434 199200 142490 200000
rect 142802 199200 142858 200000
rect 143170 199200 143226 200000
rect 143538 199200 143594 200000
rect 143906 199200 143962 200000
rect 144274 199200 144330 200000
rect 144642 199200 144698 200000
rect 145010 199200 145066 200000
rect 145378 199200 145434 200000
rect 145746 199200 145802 200000
rect 146114 199200 146170 200000
rect 146482 199200 146538 200000
rect 146850 199200 146906 200000
rect 147218 199200 147274 200000
rect 147586 199200 147642 200000
rect 147954 199200 148010 200000
rect 148322 199200 148378 200000
rect 148690 199200 148746 200000
rect 149058 199200 149114 200000
rect 149426 199200 149482 200000
rect 149794 199200 149850 200000
rect 150162 199200 150218 200000
rect 150530 199200 150586 200000
rect 150898 199200 150954 200000
rect 151266 199200 151322 200000
rect 151634 199200 151690 200000
rect 152002 199200 152058 200000
rect 152370 199200 152426 200000
rect 152738 199200 152794 200000
rect 153106 199200 153162 200000
rect 153474 199200 153530 200000
rect 153842 199200 153898 200000
rect 154210 199200 154266 200000
rect 154578 199200 154634 200000
rect 154946 199200 155002 200000
rect 155314 199200 155370 200000
rect 155682 199200 155738 200000
rect 156050 199200 156106 200000
rect 156418 199200 156474 200000
rect 156786 199200 156842 200000
rect 157154 199200 157210 200000
rect 157522 199200 157578 200000
rect 157890 199200 157946 200000
rect 158258 199200 158314 200000
rect 158626 199200 158682 200000
rect 158994 199200 159050 200000
rect 159362 199200 159418 200000
rect 159730 199200 159786 200000
rect 160098 199200 160154 200000
rect 160466 199200 160522 200000
rect 160834 199200 160890 200000
rect 161202 199200 161258 200000
rect 161570 199200 161626 200000
rect 161938 199200 161994 200000
rect 162306 199200 162362 200000
rect 162674 199200 162730 200000
rect 163042 199200 163098 200000
rect 163410 199200 163466 200000
rect 163778 199200 163834 200000
rect 164146 199200 164202 200000
rect 164514 199200 164570 200000
rect 164882 199200 164938 200000
rect 165250 199200 165306 200000
rect 165618 199200 165674 200000
rect 165986 199200 166042 200000
rect 166354 199200 166410 200000
rect 166722 199200 166778 200000
rect 167090 199200 167146 200000
rect 167458 199200 167514 200000
rect 167826 199200 167882 200000
rect 168194 199200 168250 200000
rect 168562 199200 168618 200000
rect 168930 199200 168986 200000
rect 169298 199200 169354 200000
rect 169666 199200 169722 200000
rect 170034 199200 170090 200000
rect 170402 199200 170458 200000
rect 170770 199200 170826 200000
rect 171138 199200 171194 200000
rect 171506 199200 171562 200000
rect 171874 199200 171930 200000
rect 172242 199200 172298 200000
rect 172610 199200 172666 200000
rect 172978 199200 173034 200000
rect 173346 199200 173402 200000
rect 173714 199200 173770 200000
rect 174082 199200 174138 200000
rect 174450 199200 174506 200000
rect 174818 199200 174874 200000
rect 175186 199200 175242 200000
rect 175554 199200 175610 200000
rect 175922 199200 175978 200000
rect 176290 199200 176346 200000
rect 176658 199200 176714 200000
rect 177026 199200 177082 200000
rect 177394 199200 177450 200000
rect 177762 199200 177818 200000
rect 178130 199200 178186 200000
rect 178498 199200 178554 200000
rect 178866 199200 178922 200000
rect 179234 199200 179290 200000
rect 179602 199200 179658 200000
rect 179970 199200 180026 200000
rect 180338 199200 180394 200000
rect 180706 199200 180762 200000
rect 181074 199200 181130 200000
rect 181442 199200 181498 200000
rect 181810 199200 181866 200000
rect 182178 199200 182234 200000
rect 182546 199200 182602 200000
rect 182914 199200 182970 200000
rect 183282 199200 183338 200000
rect 183650 199200 183706 200000
rect 184018 199200 184074 200000
rect 184386 199200 184442 200000
rect 184754 199200 184810 200000
rect 185122 199200 185178 200000
rect 185490 199200 185546 200000
rect 185858 199200 185914 200000
rect 186226 199200 186282 200000
rect 186594 199200 186650 200000
rect 186962 199200 187018 200000
rect 187330 199200 187386 200000
rect 187698 199200 187754 200000
rect 188066 199200 188122 200000
rect 188434 199200 188490 200000
rect 188802 199200 188858 200000
rect 189170 199200 189226 200000
rect 189538 199200 189594 200000
rect 189906 199200 189962 200000
rect 190274 199200 190330 200000
rect 190642 199200 190698 200000
rect 191010 199200 191066 200000
rect 191378 199200 191434 200000
rect 191746 199200 191802 200000
rect 192114 199200 192170 200000
rect 192482 199200 192538 200000
rect 192850 199200 192906 200000
rect 193218 199200 193274 200000
rect 193586 199200 193642 200000
rect 193954 199200 194010 200000
rect 194322 199200 194378 200000
rect 194690 199200 194746 200000
rect 195058 199200 195114 200000
rect 195426 199200 195482 200000
rect 195794 199200 195850 200000
rect 196162 199200 196218 200000
rect 1950 0 2006 800
rect 3330 0 3386 800
rect 4710 0 4766 800
rect 6090 0 6146 800
rect 7470 0 7526 800
rect 8850 0 8906 800
rect 10230 0 10286 800
rect 11610 0 11666 800
rect 12990 0 13046 800
rect 14370 0 14426 800
rect 15750 0 15806 800
rect 17130 0 17186 800
rect 18510 0 18566 800
rect 19890 0 19946 800
rect 21270 0 21326 800
rect 22650 0 22706 800
rect 24030 0 24086 800
rect 25410 0 25466 800
rect 26790 0 26846 800
rect 28170 0 28226 800
rect 29550 0 29606 800
rect 30930 0 30986 800
rect 32310 0 32366 800
rect 33690 0 33746 800
rect 35070 0 35126 800
rect 36450 0 36506 800
rect 37830 0 37886 800
rect 39210 0 39266 800
rect 40590 0 40646 800
rect 41970 0 42026 800
rect 43350 0 43406 800
rect 44730 0 44786 800
rect 46110 0 46166 800
rect 47490 0 47546 800
rect 48870 0 48926 800
rect 50250 0 50306 800
rect 51630 0 51686 800
rect 53010 0 53066 800
rect 54390 0 54446 800
rect 55770 0 55826 800
rect 57150 0 57206 800
rect 58530 0 58586 800
rect 59910 0 59966 800
rect 61290 0 61346 800
rect 62670 0 62726 800
rect 64050 0 64106 800
rect 65430 0 65486 800
rect 66810 0 66866 800
rect 68190 0 68246 800
rect 69570 0 69626 800
rect 70950 0 71006 800
rect 72330 0 72386 800
rect 73710 0 73766 800
rect 75090 0 75146 800
rect 76470 0 76526 800
rect 77850 0 77906 800
rect 79230 0 79286 800
rect 80610 0 80666 800
rect 81990 0 82046 800
rect 83370 0 83426 800
rect 84750 0 84806 800
rect 86130 0 86186 800
rect 87510 0 87566 800
rect 88890 0 88946 800
rect 90270 0 90326 800
rect 91650 0 91706 800
rect 93030 0 93086 800
rect 94410 0 94466 800
rect 95790 0 95846 800
rect 97170 0 97226 800
rect 98550 0 98606 800
rect 99930 0 99986 800
rect 101310 0 101366 800
rect 102690 0 102746 800
rect 104070 0 104126 800
rect 105450 0 105506 800
rect 106830 0 106886 800
rect 108210 0 108266 800
rect 109590 0 109646 800
rect 110970 0 111026 800
rect 112350 0 112406 800
rect 113730 0 113786 800
rect 115110 0 115166 800
rect 116490 0 116546 800
rect 117870 0 117926 800
rect 119250 0 119306 800
rect 120630 0 120686 800
rect 122010 0 122066 800
rect 123390 0 123446 800
rect 124770 0 124826 800
rect 126150 0 126206 800
rect 127530 0 127586 800
rect 128910 0 128966 800
rect 130290 0 130346 800
rect 131670 0 131726 800
rect 133050 0 133106 800
rect 134430 0 134486 800
rect 135810 0 135866 800
rect 137190 0 137246 800
rect 138570 0 138626 800
rect 139950 0 140006 800
rect 141330 0 141386 800
rect 142710 0 142766 800
rect 144090 0 144146 800
rect 145470 0 145526 800
rect 146850 0 146906 800
rect 148230 0 148286 800
rect 149610 0 149666 800
rect 150990 0 151046 800
rect 152370 0 152426 800
rect 153750 0 153806 800
rect 155130 0 155186 800
rect 156510 0 156566 800
rect 157890 0 157946 800
rect 159270 0 159326 800
rect 160650 0 160706 800
rect 162030 0 162086 800
rect 163410 0 163466 800
rect 164790 0 164846 800
rect 166170 0 166226 800
rect 167550 0 167606 800
rect 168930 0 168986 800
rect 170310 0 170366 800
rect 171690 0 171746 800
rect 173070 0 173126 800
rect 174450 0 174506 800
rect 175830 0 175886 800
rect 177210 0 177266 800
rect 178590 0 178646 800
rect 179970 0 180026 800
rect 181350 0 181406 800
rect 182730 0 182786 800
rect 184110 0 184166 800
rect 185490 0 185546 800
rect 186870 0 186926 800
rect 188250 0 188306 800
rect 189630 0 189686 800
rect 191010 0 191066 800
rect 192390 0 192446 800
rect 193770 0 193826 800
rect 195150 0 195206 800
rect 196530 0 196586 800
rect 197910 0 197966 800
<< obsm2 >>
rect 1952 199144 3642 199458
rect 3810 199144 4010 199458
rect 4178 199144 4378 199458
rect 4546 199144 4746 199458
rect 4914 199144 5114 199458
rect 5282 199144 5482 199458
rect 5650 199144 5850 199458
rect 6018 199144 6218 199458
rect 6386 199144 6586 199458
rect 6754 199144 6954 199458
rect 7122 199144 7322 199458
rect 7490 199144 7690 199458
rect 7858 199144 8058 199458
rect 8226 199144 8426 199458
rect 8594 199144 8794 199458
rect 8962 199144 9162 199458
rect 9330 199144 9530 199458
rect 9698 199144 9898 199458
rect 10066 199144 10266 199458
rect 10434 199144 10634 199458
rect 10802 199144 11002 199458
rect 11170 199144 11370 199458
rect 11538 199144 11738 199458
rect 11906 199144 12106 199458
rect 12274 199144 12474 199458
rect 12642 199144 12842 199458
rect 13010 199144 13210 199458
rect 13378 199144 13578 199458
rect 13746 199144 13946 199458
rect 14114 199144 14314 199458
rect 14482 199144 14682 199458
rect 14850 199144 15050 199458
rect 15218 199144 15418 199458
rect 15586 199144 15786 199458
rect 15954 199144 16154 199458
rect 16322 199144 16522 199458
rect 16690 199144 16890 199458
rect 17058 199144 17258 199458
rect 17426 199144 17626 199458
rect 17794 199144 17994 199458
rect 18162 199144 18362 199458
rect 18530 199144 18730 199458
rect 18898 199144 19098 199458
rect 19266 199144 19466 199458
rect 19634 199144 19834 199458
rect 20002 199144 20202 199458
rect 20370 199144 20570 199458
rect 20738 199144 20938 199458
rect 21106 199144 21306 199458
rect 21474 199144 21674 199458
rect 21842 199144 22042 199458
rect 22210 199144 22410 199458
rect 22578 199144 22778 199458
rect 22946 199144 23146 199458
rect 23314 199144 23514 199458
rect 23682 199144 23882 199458
rect 24050 199144 24250 199458
rect 24418 199144 24618 199458
rect 24786 199144 24986 199458
rect 25154 199144 25354 199458
rect 25522 199144 25722 199458
rect 25890 199144 26090 199458
rect 26258 199144 26458 199458
rect 26626 199144 26826 199458
rect 26994 199144 27194 199458
rect 27362 199144 27562 199458
rect 27730 199144 27930 199458
rect 28098 199144 28298 199458
rect 28466 199144 28666 199458
rect 28834 199144 29034 199458
rect 29202 199144 29402 199458
rect 29570 199144 29770 199458
rect 29938 199144 30138 199458
rect 30306 199144 30506 199458
rect 30674 199144 30874 199458
rect 31042 199144 31242 199458
rect 31410 199144 31610 199458
rect 31778 199144 31978 199458
rect 32146 199144 32346 199458
rect 32514 199144 32714 199458
rect 32882 199144 33082 199458
rect 33250 199144 33450 199458
rect 33618 199144 33818 199458
rect 33986 199144 34186 199458
rect 34354 199144 34554 199458
rect 34722 199144 34922 199458
rect 35090 199144 35290 199458
rect 35458 199144 35658 199458
rect 35826 199144 36026 199458
rect 36194 199144 36394 199458
rect 36562 199144 36762 199458
rect 36930 199144 37130 199458
rect 37298 199144 37498 199458
rect 37666 199144 37866 199458
rect 38034 199144 38234 199458
rect 38402 199144 38602 199458
rect 38770 199144 38970 199458
rect 39138 199144 39338 199458
rect 39506 199144 39706 199458
rect 39874 199144 40074 199458
rect 40242 199144 40442 199458
rect 40610 199144 40810 199458
rect 40978 199144 41178 199458
rect 41346 199144 41546 199458
rect 41714 199144 41914 199458
rect 42082 199144 42282 199458
rect 42450 199144 42650 199458
rect 42818 199144 43018 199458
rect 43186 199144 43386 199458
rect 43554 199144 43754 199458
rect 43922 199144 44122 199458
rect 44290 199144 44490 199458
rect 44658 199144 44858 199458
rect 45026 199144 45226 199458
rect 45394 199144 45594 199458
rect 45762 199144 45962 199458
rect 46130 199144 46330 199458
rect 46498 199144 46698 199458
rect 46866 199144 47066 199458
rect 47234 199144 47434 199458
rect 47602 199144 47802 199458
rect 47970 199144 48170 199458
rect 48338 199144 48538 199458
rect 48706 199144 48906 199458
rect 49074 199144 49274 199458
rect 49442 199144 49642 199458
rect 49810 199144 50010 199458
rect 50178 199144 50378 199458
rect 50546 199144 50746 199458
rect 50914 199144 51114 199458
rect 51282 199144 51482 199458
rect 51650 199144 51850 199458
rect 52018 199144 52218 199458
rect 52386 199144 52586 199458
rect 52754 199144 52954 199458
rect 53122 199144 53322 199458
rect 53490 199144 53690 199458
rect 53858 199144 54058 199458
rect 54226 199144 54426 199458
rect 54594 199144 54794 199458
rect 54962 199144 55162 199458
rect 55330 199144 55530 199458
rect 55698 199144 55898 199458
rect 56066 199144 56266 199458
rect 56434 199144 56634 199458
rect 56802 199144 57002 199458
rect 57170 199144 57370 199458
rect 57538 199144 57738 199458
rect 57906 199144 58106 199458
rect 58274 199144 58474 199458
rect 58642 199144 58842 199458
rect 59010 199144 59210 199458
rect 59378 199144 59578 199458
rect 59746 199144 59946 199458
rect 60114 199144 60314 199458
rect 60482 199144 60682 199458
rect 60850 199144 61050 199458
rect 61218 199144 61418 199458
rect 61586 199144 61786 199458
rect 61954 199144 62154 199458
rect 62322 199144 62522 199458
rect 62690 199144 62890 199458
rect 63058 199144 63258 199458
rect 63426 199144 63626 199458
rect 63794 199144 63994 199458
rect 64162 199144 64362 199458
rect 64530 199144 64730 199458
rect 64898 199144 65098 199458
rect 65266 199144 65466 199458
rect 65634 199144 65834 199458
rect 66002 199144 66202 199458
rect 66370 199144 66570 199458
rect 66738 199144 66938 199458
rect 67106 199144 67306 199458
rect 67474 199144 67674 199458
rect 67842 199144 68042 199458
rect 68210 199144 68410 199458
rect 68578 199144 68778 199458
rect 68946 199144 69146 199458
rect 69314 199144 69514 199458
rect 69682 199144 69882 199458
rect 70050 199144 70250 199458
rect 70418 199144 70618 199458
rect 70786 199144 70986 199458
rect 71154 199144 71354 199458
rect 71522 199144 71722 199458
rect 71890 199144 72090 199458
rect 72258 199144 72458 199458
rect 72626 199144 72826 199458
rect 72994 199144 73194 199458
rect 73362 199144 73562 199458
rect 73730 199144 73930 199458
rect 74098 199144 74298 199458
rect 74466 199144 74666 199458
rect 74834 199144 75034 199458
rect 75202 199144 75402 199458
rect 75570 199144 75770 199458
rect 75938 199144 76138 199458
rect 76306 199144 76506 199458
rect 76674 199144 76874 199458
rect 77042 199144 77242 199458
rect 77410 199144 77610 199458
rect 77778 199144 77978 199458
rect 78146 199144 78346 199458
rect 78514 199144 78714 199458
rect 78882 199144 79082 199458
rect 79250 199144 79450 199458
rect 79618 199144 79818 199458
rect 79986 199144 80186 199458
rect 80354 199144 80554 199458
rect 80722 199144 80922 199458
rect 81090 199144 81290 199458
rect 81458 199144 81658 199458
rect 81826 199144 82026 199458
rect 82194 199144 82394 199458
rect 82562 199144 82762 199458
rect 82930 199144 83130 199458
rect 83298 199144 83498 199458
rect 83666 199144 83866 199458
rect 84034 199144 84234 199458
rect 84402 199144 84602 199458
rect 84770 199144 84970 199458
rect 85138 199144 85338 199458
rect 85506 199144 85706 199458
rect 85874 199144 86074 199458
rect 86242 199144 86442 199458
rect 86610 199144 86810 199458
rect 86978 199144 87178 199458
rect 87346 199144 87546 199458
rect 87714 199144 87914 199458
rect 88082 199144 88282 199458
rect 88450 199144 88650 199458
rect 88818 199144 89018 199458
rect 89186 199144 89386 199458
rect 89554 199144 89754 199458
rect 89922 199144 90122 199458
rect 90290 199144 90490 199458
rect 90658 199144 90858 199458
rect 91026 199144 91226 199458
rect 91394 199144 91594 199458
rect 91762 199144 91962 199458
rect 92130 199144 92330 199458
rect 92498 199144 92698 199458
rect 92866 199144 93066 199458
rect 93234 199144 93434 199458
rect 93602 199144 93802 199458
rect 93970 199144 94170 199458
rect 94338 199144 94538 199458
rect 94706 199144 94906 199458
rect 95074 199144 95274 199458
rect 95442 199144 95642 199458
rect 95810 199144 96010 199458
rect 96178 199144 96378 199458
rect 96546 199144 96746 199458
rect 96914 199144 97114 199458
rect 97282 199144 97482 199458
rect 97650 199144 97850 199458
rect 98018 199144 98218 199458
rect 98386 199144 98586 199458
rect 98754 199144 98954 199458
rect 99122 199144 99322 199458
rect 99490 199144 99690 199458
rect 99858 199144 100058 199458
rect 100226 199144 100426 199458
rect 100594 199144 100794 199458
rect 100962 199144 101162 199458
rect 101330 199144 101530 199458
rect 101698 199144 101898 199458
rect 102066 199144 102266 199458
rect 102434 199144 102634 199458
rect 102802 199144 103002 199458
rect 103170 199144 103370 199458
rect 103538 199144 103738 199458
rect 103906 199144 104106 199458
rect 104274 199144 104474 199458
rect 104642 199144 104842 199458
rect 105010 199144 105210 199458
rect 105378 199144 105578 199458
rect 105746 199144 105946 199458
rect 106114 199144 106314 199458
rect 106482 199144 106682 199458
rect 106850 199144 107050 199458
rect 107218 199144 107418 199458
rect 107586 199144 107786 199458
rect 107954 199144 108154 199458
rect 108322 199144 108522 199458
rect 108690 199144 108890 199458
rect 109058 199144 109258 199458
rect 109426 199144 109626 199458
rect 109794 199144 109994 199458
rect 110162 199144 110362 199458
rect 110530 199144 110730 199458
rect 110898 199144 111098 199458
rect 111266 199144 111466 199458
rect 111634 199144 111834 199458
rect 112002 199144 112202 199458
rect 112370 199144 112570 199458
rect 112738 199144 112938 199458
rect 113106 199144 113306 199458
rect 113474 199144 113674 199458
rect 113842 199144 114042 199458
rect 114210 199144 114410 199458
rect 114578 199144 114778 199458
rect 114946 199144 115146 199458
rect 115314 199144 115514 199458
rect 115682 199144 115882 199458
rect 116050 199144 116250 199458
rect 116418 199144 116618 199458
rect 116786 199144 116986 199458
rect 117154 199144 117354 199458
rect 117522 199144 117722 199458
rect 117890 199144 118090 199458
rect 118258 199144 118458 199458
rect 118626 199144 118826 199458
rect 118994 199144 119194 199458
rect 119362 199144 119562 199458
rect 119730 199144 119930 199458
rect 120098 199144 120298 199458
rect 120466 199144 120666 199458
rect 120834 199144 121034 199458
rect 121202 199144 121402 199458
rect 121570 199144 121770 199458
rect 121938 199144 122138 199458
rect 122306 199144 122506 199458
rect 122674 199144 122874 199458
rect 123042 199144 123242 199458
rect 123410 199144 123610 199458
rect 123778 199144 123978 199458
rect 124146 199144 124346 199458
rect 124514 199144 124714 199458
rect 124882 199144 125082 199458
rect 125250 199144 125450 199458
rect 125618 199144 125818 199458
rect 125986 199144 126186 199458
rect 126354 199144 126554 199458
rect 126722 199144 126922 199458
rect 127090 199144 127290 199458
rect 127458 199144 127658 199458
rect 127826 199144 128026 199458
rect 128194 199144 128394 199458
rect 128562 199144 128762 199458
rect 128930 199144 129130 199458
rect 129298 199144 129498 199458
rect 129666 199144 129866 199458
rect 130034 199144 130234 199458
rect 130402 199144 130602 199458
rect 130770 199144 130970 199458
rect 131138 199144 131338 199458
rect 131506 199144 131706 199458
rect 131874 199144 132074 199458
rect 132242 199144 132442 199458
rect 132610 199144 132810 199458
rect 132978 199144 133178 199458
rect 133346 199144 133546 199458
rect 133714 199144 133914 199458
rect 134082 199144 134282 199458
rect 134450 199144 134650 199458
rect 134818 199144 135018 199458
rect 135186 199144 135386 199458
rect 135554 199144 135754 199458
rect 135922 199144 136122 199458
rect 136290 199144 136490 199458
rect 136658 199144 136858 199458
rect 137026 199144 137226 199458
rect 137394 199144 137594 199458
rect 137762 199144 137962 199458
rect 138130 199144 138330 199458
rect 138498 199144 138698 199458
rect 138866 199144 139066 199458
rect 139234 199144 139434 199458
rect 139602 199144 139802 199458
rect 139970 199144 140170 199458
rect 140338 199144 140538 199458
rect 140706 199144 140906 199458
rect 141074 199144 141274 199458
rect 141442 199144 141642 199458
rect 141810 199144 142010 199458
rect 142178 199144 142378 199458
rect 142546 199144 142746 199458
rect 142914 199144 143114 199458
rect 143282 199144 143482 199458
rect 143650 199144 143850 199458
rect 144018 199144 144218 199458
rect 144386 199144 144586 199458
rect 144754 199144 144954 199458
rect 145122 199144 145322 199458
rect 145490 199144 145690 199458
rect 145858 199144 146058 199458
rect 146226 199144 146426 199458
rect 146594 199144 146794 199458
rect 146962 199144 147162 199458
rect 147330 199144 147530 199458
rect 147698 199144 147898 199458
rect 148066 199144 148266 199458
rect 148434 199144 148634 199458
rect 148802 199144 149002 199458
rect 149170 199144 149370 199458
rect 149538 199144 149738 199458
rect 149906 199144 150106 199458
rect 150274 199144 150474 199458
rect 150642 199144 150842 199458
rect 151010 199144 151210 199458
rect 151378 199144 151578 199458
rect 151746 199144 151946 199458
rect 152114 199144 152314 199458
rect 152482 199144 152682 199458
rect 152850 199144 153050 199458
rect 153218 199144 153418 199458
rect 153586 199144 153786 199458
rect 153954 199144 154154 199458
rect 154322 199144 154522 199458
rect 154690 199144 154890 199458
rect 155058 199144 155258 199458
rect 155426 199144 155626 199458
rect 155794 199144 155994 199458
rect 156162 199144 156362 199458
rect 156530 199144 156730 199458
rect 156898 199144 157098 199458
rect 157266 199144 157466 199458
rect 157634 199144 157834 199458
rect 158002 199144 158202 199458
rect 158370 199144 158570 199458
rect 158738 199144 158938 199458
rect 159106 199144 159306 199458
rect 159474 199144 159674 199458
rect 159842 199144 160042 199458
rect 160210 199144 160410 199458
rect 160578 199144 160778 199458
rect 160946 199144 161146 199458
rect 161314 199144 161514 199458
rect 161682 199144 161882 199458
rect 162050 199144 162250 199458
rect 162418 199144 162618 199458
rect 162786 199144 162986 199458
rect 163154 199144 163354 199458
rect 163522 199144 163722 199458
rect 163890 199144 164090 199458
rect 164258 199144 164458 199458
rect 164626 199144 164826 199458
rect 164994 199144 165194 199458
rect 165362 199144 165562 199458
rect 165730 199144 165930 199458
rect 166098 199144 166298 199458
rect 166466 199144 166666 199458
rect 166834 199144 167034 199458
rect 167202 199144 167402 199458
rect 167570 199144 167770 199458
rect 167938 199144 168138 199458
rect 168306 199144 168506 199458
rect 168674 199144 168874 199458
rect 169042 199144 169242 199458
rect 169410 199144 169610 199458
rect 169778 199144 169978 199458
rect 170146 199144 170346 199458
rect 170514 199144 170714 199458
rect 170882 199144 171082 199458
rect 171250 199144 171450 199458
rect 171618 199144 171818 199458
rect 171986 199144 172186 199458
rect 172354 199144 172554 199458
rect 172722 199144 172922 199458
rect 173090 199144 173290 199458
rect 173458 199144 173658 199458
rect 173826 199144 174026 199458
rect 174194 199144 174394 199458
rect 174562 199144 174762 199458
rect 174930 199144 175130 199458
rect 175298 199144 175498 199458
rect 175666 199144 175866 199458
rect 176034 199144 176234 199458
rect 176402 199144 176602 199458
rect 176770 199144 176970 199458
rect 177138 199144 177338 199458
rect 177506 199144 177706 199458
rect 177874 199144 178074 199458
rect 178242 199144 178442 199458
rect 178610 199144 178810 199458
rect 178978 199144 179178 199458
rect 179346 199144 179546 199458
rect 179714 199144 179914 199458
rect 180082 199144 180282 199458
rect 180450 199144 180650 199458
rect 180818 199144 181018 199458
rect 181186 199144 181386 199458
rect 181554 199144 181754 199458
rect 181922 199144 182122 199458
rect 182290 199144 182490 199458
rect 182658 199144 182858 199458
rect 183026 199144 183226 199458
rect 183394 199144 183594 199458
rect 183762 199144 183962 199458
rect 184130 199144 184330 199458
rect 184498 199144 184698 199458
rect 184866 199144 185066 199458
rect 185234 199144 185434 199458
rect 185602 199144 185802 199458
rect 185970 199144 186170 199458
rect 186338 199144 186538 199458
rect 186706 199144 186906 199458
rect 187074 199144 187274 199458
rect 187442 199144 187642 199458
rect 187810 199144 188010 199458
rect 188178 199144 188378 199458
rect 188546 199144 188746 199458
rect 188914 199144 189114 199458
rect 189282 199144 189482 199458
rect 189650 199144 189850 199458
rect 190018 199144 190218 199458
rect 190386 199144 190586 199458
rect 190754 199144 190954 199458
rect 191122 199144 191322 199458
rect 191490 199144 191690 199458
rect 191858 199144 192058 199458
rect 192226 199144 192426 199458
rect 192594 199144 192794 199458
rect 192962 199144 193162 199458
rect 193330 199144 193530 199458
rect 193698 199144 193898 199458
rect 194066 199144 194266 199458
rect 194434 199144 194634 199458
rect 194802 199144 195002 199458
rect 195170 199144 195370 199458
rect 195538 199144 195738 199458
rect 195906 199144 196106 199458
rect 196274 199144 197964 199458
rect 1952 856 197964 199144
rect 2062 734 3274 856
rect 3442 734 4654 856
rect 4822 734 6034 856
rect 6202 734 7414 856
rect 7582 734 8794 856
rect 8962 734 10174 856
rect 10342 734 11554 856
rect 11722 734 12934 856
rect 13102 734 14314 856
rect 14482 734 15694 856
rect 15862 734 17074 856
rect 17242 734 18454 856
rect 18622 734 19834 856
rect 20002 734 21214 856
rect 21382 734 22594 856
rect 22762 734 23974 856
rect 24142 734 25354 856
rect 25522 734 26734 856
rect 26902 734 28114 856
rect 28282 734 29494 856
rect 29662 734 30874 856
rect 31042 734 32254 856
rect 32422 734 33634 856
rect 33802 734 35014 856
rect 35182 734 36394 856
rect 36562 734 37774 856
rect 37942 734 39154 856
rect 39322 734 40534 856
rect 40702 734 41914 856
rect 42082 734 43294 856
rect 43462 734 44674 856
rect 44842 734 46054 856
rect 46222 734 47434 856
rect 47602 734 48814 856
rect 48982 734 50194 856
rect 50362 734 51574 856
rect 51742 734 52954 856
rect 53122 734 54334 856
rect 54502 734 55714 856
rect 55882 734 57094 856
rect 57262 734 58474 856
rect 58642 734 59854 856
rect 60022 734 61234 856
rect 61402 734 62614 856
rect 62782 734 63994 856
rect 64162 734 65374 856
rect 65542 734 66754 856
rect 66922 734 68134 856
rect 68302 734 69514 856
rect 69682 734 70894 856
rect 71062 734 72274 856
rect 72442 734 73654 856
rect 73822 734 75034 856
rect 75202 734 76414 856
rect 76582 734 77794 856
rect 77962 734 79174 856
rect 79342 734 80554 856
rect 80722 734 81934 856
rect 82102 734 83314 856
rect 83482 734 84694 856
rect 84862 734 86074 856
rect 86242 734 87454 856
rect 87622 734 88834 856
rect 89002 734 90214 856
rect 90382 734 91594 856
rect 91762 734 92974 856
rect 93142 734 94354 856
rect 94522 734 95734 856
rect 95902 734 97114 856
rect 97282 734 98494 856
rect 98662 734 99874 856
rect 100042 734 101254 856
rect 101422 734 102634 856
rect 102802 734 104014 856
rect 104182 734 105394 856
rect 105562 734 106774 856
rect 106942 734 108154 856
rect 108322 734 109534 856
rect 109702 734 110914 856
rect 111082 734 112294 856
rect 112462 734 113674 856
rect 113842 734 115054 856
rect 115222 734 116434 856
rect 116602 734 117814 856
rect 117982 734 119194 856
rect 119362 734 120574 856
rect 120742 734 121954 856
rect 122122 734 123334 856
rect 123502 734 124714 856
rect 124882 734 126094 856
rect 126262 734 127474 856
rect 127642 734 128854 856
rect 129022 734 130234 856
rect 130402 734 131614 856
rect 131782 734 132994 856
rect 133162 734 134374 856
rect 134542 734 135754 856
rect 135922 734 137134 856
rect 137302 734 138514 856
rect 138682 734 139894 856
rect 140062 734 141274 856
rect 141442 734 142654 856
rect 142822 734 144034 856
rect 144202 734 145414 856
rect 145582 734 146794 856
rect 146962 734 148174 856
rect 148342 734 149554 856
rect 149722 734 150934 856
rect 151102 734 152314 856
rect 152482 734 153694 856
rect 153862 734 155074 856
rect 155242 734 156454 856
rect 156622 734 157834 856
rect 158002 734 159214 856
rect 159382 734 160594 856
rect 160762 734 161974 856
rect 162142 734 163354 856
rect 163522 734 164734 856
rect 164902 734 166114 856
rect 166282 734 167494 856
rect 167662 734 168874 856
rect 169042 734 170254 856
rect 170422 734 171634 856
rect 171802 734 173014 856
rect 173182 734 174394 856
rect 174562 734 175774 856
rect 175942 734 177154 856
rect 177322 734 178534 856
rect 178702 734 179914 856
rect 180082 734 181294 856
rect 181462 734 182674 856
rect 182842 734 184054 856
rect 184222 734 185434 856
rect 185602 734 186814 856
rect 186982 734 188194 856
rect 188362 734 189574 856
rect 189742 734 190954 856
rect 191122 734 192334 856
rect 192502 734 193714 856
rect 193882 734 195094 856
rect 195262 734 196474 856
rect 196642 734 197854 856
<< obsm3 >>
rect 4210 1803 197511 199476
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
<< obsm4 >>
rect 68139 197600 174005 199477
rect 68139 2048 80928 197600
rect 81408 2048 96288 197600
rect 96768 2048 111648 197600
rect 112128 2048 127008 197600
rect 127488 2048 142368 197600
rect 142848 2048 157728 197600
rect 158208 2048 173088 197600
rect 173568 2048 174005 197600
rect 68139 1803 174005 2048
<< labels >>
rlabel metal2 s 193770 0 193826 800 6 Serial_input
port 1 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 Serial_output
port 2 nsew signal output
rlabel metal2 s 188250 0 188306 800 6 clk
port 3 nsew signal output
rlabel metal2 s 71778 199200 71834 200000 6 data_mem_addr[0]
port 4 nsew signal output
rlabel metal2 s 73250 199200 73306 200000 6 data_mem_addr[1]
port 5 nsew signal output
rlabel metal2 s 74722 199200 74778 200000 6 data_mem_addr[2]
port 6 nsew signal output
rlabel metal2 s 76194 199200 76250 200000 6 data_mem_addr[3]
port 7 nsew signal output
rlabel metal2 s 77666 199200 77722 200000 6 data_mem_addr[4]
port 8 nsew signal output
rlabel metal2 s 78770 199200 78826 200000 6 data_mem_addr[5]
port 9 nsew signal output
rlabel metal2 s 79874 199200 79930 200000 6 data_mem_addr[6]
port 10 nsew signal output
rlabel metal2 s 80978 199200 81034 200000 6 data_mem_addr[7]
port 11 nsew signal output
rlabel metal2 s 71410 199200 71466 200000 6 data_mem_csb
port 12 nsew signal output
rlabel metal2 s 72146 199200 72202 200000 6 data_read_data[0]
port 13 nsew signal input
rlabel metal2 s 83554 199200 83610 200000 6 data_read_data[10]
port 14 nsew signal input
rlabel metal2 s 84290 199200 84346 200000 6 data_read_data[11]
port 15 nsew signal input
rlabel metal2 s 85026 199200 85082 200000 6 data_read_data[12]
port 16 nsew signal input
rlabel metal2 s 85762 199200 85818 200000 6 data_read_data[13]
port 17 nsew signal input
rlabel metal2 s 86498 199200 86554 200000 6 data_read_data[14]
port 18 nsew signal input
rlabel metal2 s 87234 199200 87290 200000 6 data_read_data[15]
port 19 nsew signal input
rlabel metal2 s 73618 199200 73674 200000 6 data_read_data[1]
port 20 nsew signal input
rlabel metal2 s 75090 199200 75146 200000 6 data_read_data[2]
port 21 nsew signal input
rlabel metal2 s 76562 199200 76618 200000 6 data_read_data[3]
port 22 nsew signal input
rlabel metal2 s 78034 199200 78090 200000 6 data_read_data[4]
port 23 nsew signal input
rlabel metal2 s 79138 199200 79194 200000 6 data_read_data[5]
port 24 nsew signal input
rlabel metal2 s 80242 199200 80298 200000 6 data_read_data[6]
port 25 nsew signal input
rlabel metal2 s 81346 199200 81402 200000 6 data_read_data[7]
port 26 nsew signal input
rlabel metal2 s 82082 199200 82138 200000 6 data_read_data[8]
port 27 nsew signal input
rlabel metal2 s 82818 199200 82874 200000 6 data_read_data[9]
port 28 nsew signal input
rlabel metal2 s 72514 199200 72570 200000 6 data_wmask[0]
port 29 nsew signal output
rlabel metal2 s 73986 199200 74042 200000 6 data_wmask[1]
port 30 nsew signal output
rlabel metal2 s 75458 199200 75514 200000 6 data_wmask[2]
port 31 nsew signal output
rlabel metal2 s 76930 199200 76986 200000 6 data_wmask[3]
port 32 nsew signal output
rlabel metal2 s 72882 199200 72938 200000 6 data_write_data[0]
port 33 nsew signal output
rlabel metal2 s 83922 199200 83978 200000 6 data_write_data[10]
port 34 nsew signal output
rlabel metal2 s 84658 199200 84714 200000 6 data_write_data[11]
port 35 nsew signal output
rlabel metal2 s 85394 199200 85450 200000 6 data_write_data[12]
port 36 nsew signal output
rlabel metal2 s 86130 199200 86186 200000 6 data_write_data[13]
port 37 nsew signal output
rlabel metal2 s 86866 199200 86922 200000 6 data_write_data[14]
port 38 nsew signal output
rlabel metal2 s 87602 199200 87658 200000 6 data_write_data[15]
port 39 nsew signal output
rlabel metal2 s 74354 199200 74410 200000 6 data_write_data[1]
port 40 nsew signal output
rlabel metal2 s 75826 199200 75882 200000 6 data_write_data[2]
port 41 nsew signal output
rlabel metal2 s 77298 199200 77354 200000 6 data_write_data[3]
port 42 nsew signal output
rlabel metal2 s 78402 199200 78458 200000 6 data_write_data[4]
port 43 nsew signal output
rlabel metal2 s 79506 199200 79562 200000 6 data_write_data[5]
port 44 nsew signal output
rlabel metal2 s 80610 199200 80666 200000 6 data_write_data[6]
port 45 nsew signal output
rlabel metal2 s 81714 199200 81770 200000 6 data_write_data[7]
port 46 nsew signal output
rlabel metal2 s 82450 199200 82506 200000 6 data_write_data[8]
port 47 nsew signal output
rlabel metal2 s 83186 199200 83242 200000 6 data_write_data[9]
port 48 nsew signal output
rlabel metal2 s 87970 199200 88026 200000 6 dataw_enb
port 49 nsew signal output
rlabel metal2 s 196530 0 196586 800 6 high
port 50 nsew signal output
rlabel metal2 s 192390 0 192446 800 6 hlt
port 51 nsew signal input
rlabel metal2 s 88338 199200 88394 200000 6 instr_mem_addr_9bit[0]
port 52 nsew signal output
rlabel metal2 s 92754 199200 92810 200000 6 instr_mem_addr_9bit[1]
port 53 nsew signal output
rlabel metal2 s 97170 199200 97226 200000 6 instr_mem_addr_9bit[2]
port 54 nsew signal output
rlabel metal2 s 101586 199200 101642 200000 6 instr_mem_addr_9bit[3]
port 55 nsew signal output
rlabel metal2 s 106002 199200 106058 200000 6 instr_mem_addr_9bit[4]
port 56 nsew signal output
rlabel metal2 s 110050 199200 110106 200000 6 instr_mem_addr_9bit[5]
port 57 nsew signal output
rlabel metal2 s 114098 199200 114154 200000 6 instr_mem_addr_9bit[6]
port 58 nsew signal output
rlabel metal2 s 118146 199200 118202 200000 6 instr_mem_addr_9bit[7]
port 59 nsew signal output
rlabel metal2 s 122194 199200 122250 200000 6 instr_mem_addr_9bit[8]
port 60 nsew signal output
rlabel metal2 s 88706 199200 88762 200000 6 instr_mem_csb[0]
port 61 nsew signal output
rlabel metal2 s 93122 199200 93178 200000 6 instr_mem_csb[1]
port 62 nsew signal output
rlabel metal2 s 97538 199200 97594 200000 6 instr_mem_csb[2]
port 63 nsew signal output
rlabel metal2 s 101954 199200 102010 200000 6 instr_mem_csb[3]
port 64 nsew signal output
rlabel metal2 s 106370 199200 106426 200000 6 instr_mem_csb[4]
port 65 nsew signal output
rlabel metal2 s 110418 199200 110474 200000 6 instr_mem_csb[5]
port 66 nsew signal output
rlabel metal2 s 114466 199200 114522 200000 6 instr_mem_csb[6]
port 67 nsew signal output
rlabel metal2 s 118514 199200 118570 200000 6 instr_mem_csb[7]
port 68 nsew signal output
rlabel metal2 s 89074 199200 89130 200000 6 instr_read_data0[0]
port 69 nsew signal input
rlabel metal2 s 129186 199200 129242 200000 6 instr_read_data0[10]
port 70 nsew signal input
rlabel metal2 s 132498 199200 132554 200000 6 instr_read_data0[11]
port 71 nsew signal input
rlabel metal2 s 135810 199200 135866 200000 6 instr_read_data0[12]
port 72 nsew signal input
rlabel metal2 s 139122 199200 139178 200000 6 instr_read_data0[13]
port 73 nsew signal input
rlabel metal2 s 142434 199200 142490 200000 6 instr_read_data0[14]
port 74 nsew signal input
rlabel metal2 s 145746 199200 145802 200000 6 instr_read_data0[15]
port 75 nsew signal input
rlabel metal2 s 149058 199200 149114 200000 6 instr_read_data0[16]
port 76 nsew signal input
rlabel metal2 s 152002 199200 152058 200000 6 instr_read_data0[17]
port 77 nsew signal input
rlabel metal2 s 154946 199200 155002 200000 6 instr_read_data0[18]
port 78 nsew signal input
rlabel metal2 s 157890 199200 157946 200000 6 instr_read_data0[19]
port 79 nsew signal input
rlabel metal2 s 93490 199200 93546 200000 6 instr_read_data0[1]
port 80 nsew signal input
rlabel metal2 s 160834 199200 160890 200000 6 instr_read_data0[20]
port 81 nsew signal input
rlabel metal2 s 163778 199200 163834 200000 6 instr_read_data0[21]
port 82 nsew signal input
rlabel metal2 s 166722 199200 166778 200000 6 instr_read_data0[22]
port 83 nsew signal input
rlabel metal2 s 169666 199200 169722 200000 6 instr_read_data0[23]
port 84 nsew signal input
rlabel metal2 s 172610 199200 172666 200000 6 instr_read_data0[24]
port 85 nsew signal input
rlabel metal2 s 175554 199200 175610 200000 6 instr_read_data0[25]
port 86 nsew signal input
rlabel metal2 s 178498 199200 178554 200000 6 instr_read_data0[26]
port 87 nsew signal input
rlabel metal2 s 181442 199200 181498 200000 6 instr_read_data0[27]
port 88 nsew signal input
rlabel metal2 s 184386 199200 184442 200000 6 instr_read_data0[28]
port 89 nsew signal input
rlabel metal2 s 187330 199200 187386 200000 6 instr_read_data0[29]
port 90 nsew signal input
rlabel metal2 s 97906 199200 97962 200000 6 instr_read_data0[2]
port 91 nsew signal input
rlabel metal2 s 190274 199200 190330 200000 6 instr_read_data0[30]
port 92 nsew signal input
rlabel metal2 s 193218 199200 193274 200000 6 instr_read_data0[31]
port 93 nsew signal input
rlabel metal2 s 102322 199200 102378 200000 6 instr_read_data0[3]
port 94 nsew signal input
rlabel metal2 s 106738 199200 106794 200000 6 instr_read_data0[4]
port 95 nsew signal input
rlabel metal2 s 110786 199200 110842 200000 6 instr_read_data0[5]
port 96 nsew signal input
rlabel metal2 s 114834 199200 114890 200000 6 instr_read_data0[6]
port 97 nsew signal input
rlabel metal2 s 118882 199200 118938 200000 6 instr_read_data0[7]
port 98 nsew signal input
rlabel metal2 s 122562 199200 122618 200000 6 instr_read_data0[8]
port 99 nsew signal input
rlabel metal2 s 125874 199200 125930 200000 6 instr_read_data0[9]
port 100 nsew signal input
rlabel metal2 s 89442 199200 89498 200000 6 instr_read_data1[0]
port 101 nsew signal input
rlabel metal2 s 129554 199200 129610 200000 6 instr_read_data1[10]
port 102 nsew signal input
rlabel metal2 s 132866 199200 132922 200000 6 instr_read_data1[11]
port 103 nsew signal input
rlabel metal2 s 136178 199200 136234 200000 6 instr_read_data1[12]
port 104 nsew signal input
rlabel metal2 s 139490 199200 139546 200000 6 instr_read_data1[13]
port 105 nsew signal input
rlabel metal2 s 142802 199200 142858 200000 6 instr_read_data1[14]
port 106 nsew signal input
rlabel metal2 s 146114 199200 146170 200000 6 instr_read_data1[15]
port 107 nsew signal input
rlabel metal2 s 149426 199200 149482 200000 6 instr_read_data1[16]
port 108 nsew signal input
rlabel metal2 s 152370 199200 152426 200000 6 instr_read_data1[17]
port 109 nsew signal input
rlabel metal2 s 155314 199200 155370 200000 6 instr_read_data1[18]
port 110 nsew signal input
rlabel metal2 s 158258 199200 158314 200000 6 instr_read_data1[19]
port 111 nsew signal input
rlabel metal2 s 93858 199200 93914 200000 6 instr_read_data1[1]
port 112 nsew signal input
rlabel metal2 s 161202 199200 161258 200000 6 instr_read_data1[20]
port 113 nsew signal input
rlabel metal2 s 164146 199200 164202 200000 6 instr_read_data1[21]
port 114 nsew signal input
rlabel metal2 s 167090 199200 167146 200000 6 instr_read_data1[22]
port 115 nsew signal input
rlabel metal2 s 170034 199200 170090 200000 6 instr_read_data1[23]
port 116 nsew signal input
rlabel metal2 s 172978 199200 173034 200000 6 instr_read_data1[24]
port 117 nsew signal input
rlabel metal2 s 175922 199200 175978 200000 6 instr_read_data1[25]
port 118 nsew signal input
rlabel metal2 s 178866 199200 178922 200000 6 instr_read_data1[26]
port 119 nsew signal input
rlabel metal2 s 181810 199200 181866 200000 6 instr_read_data1[27]
port 120 nsew signal input
rlabel metal2 s 184754 199200 184810 200000 6 instr_read_data1[28]
port 121 nsew signal input
rlabel metal2 s 187698 199200 187754 200000 6 instr_read_data1[29]
port 122 nsew signal input
rlabel metal2 s 98274 199200 98330 200000 6 instr_read_data1[2]
port 123 nsew signal input
rlabel metal2 s 190642 199200 190698 200000 6 instr_read_data1[30]
port 124 nsew signal input
rlabel metal2 s 193586 199200 193642 200000 6 instr_read_data1[31]
port 125 nsew signal input
rlabel metal2 s 102690 199200 102746 200000 6 instr_read_data1[3]
port 126 nsew signal input
rlabel metal2 s 107106 199200 107162 200000 6 instr_read_data1[4]
port 127 nsew signal input
rlabel metal2 s 111154 199200 111210 200000 6 instr_read_data1[5]
port 128 nsew signal input
rlabel metal2 s 115202 199200 115258 200000 6 instr_read_data1[6]
port 129 nsew signal input
rlabel metal2 s 119250 199200 119306 200000 6 instr_read_data1[7]
port 130 nsew signal input
rlabel metal2 s 122930 199200 122986 200000 6 instr_read_data1[8]
port 131 nsew signal input
rlabel metal2 s 126242 199200 126298 200000 6 instr_read_data1[9]
port 132 nsew signal input
rlabel metal2 s 89810 199200 89866 200000 6 instr_read_data2[0]
port 133 nsew signal input
rlabel metal2 s 129922 199200 129978 200000 6 instr_read_data2[10]
port 134 nsew signal input
rlabel metal2 s 133234 199200 133290 200000 6 instr_read_data2[11]
port 135 nsew signal input
rlabel metal2 s 136546 199200 136602 200000 6 instr_read_data2[12]
port 136 nsew signal input
rlabel metal2 s 139858 199200 139914 200000 6 instr_read_data2[13]
port 137 nsew signal input
rlabel metal2 s 143170 199200 143226 200000 6 instr_read_data2[14]
port 138 nsew signal input
rlabel metal2 s 146482 199200 146538 200000 6 instr_read_data2[15]
port 139 nsew signal input
rlabel metal2 s 149794 199200 149850 200000 6 instr_read_data2[16]
port 140 nsew signal input
rlabel metal2 s 152738 199200 152794 200000 6 instr_read_data2[17]
port 141 nsew signal input
rlabel metal2 s 155682 199200 155738 200000 6 instr_read_data2[18]
port 142 nsew signal input
rlabel metal2 s 158626 199200 158682 200000 6 instr_read_data2[19]
port 143 nsew signal input
rlabel metal2 s 94226 199200 94282 200000 6 instr_read_data2[1]
port 144 nsew signal input
rlabel metal2 s 161570 199200 161626 200000 6 instr_read_data2[20]
port 145 nsew signal input
rlabel metal2 s 164514 199200 164570 200000 6 instr_read_data2[21]
port 146 nsew signal input
rlabel metal2 s 167458 199200 167514 200000 6 instr_read_data2[22]
port 147 nsew signal input
rlabel metal2 s 170402 199200 170458 200000 6 instr_read_data2[23]
port 148 nsew signal input
rlabel metal2 s 173346 199200 173402 200000 6 instr_read_data2[24]
port 149 nsew signal input
rlabel metal2 s 176290 199200 176346 200000 6 instr_read_data2[25]
port 150 nsew signal input
rlabel metal2 s 179234 199200 179290 200000 6 instr_read_data2[26]
port 151 nsew signal input
rlabel metal2 s 182178 199200 182234 200000 6 instr_read_data2[27]
port 152 nsew signal input
rlabel metal2 s 185122 199200 185178 200000 6 instr_read_data2[28]
port 153 nsew signal input
rlabel metal2 s 188066 199200 188122 200000 6 instr_read_data2[29]
port 154 nsew signal input
rlabel metal2 s 98642 199200 98698 200000 6 instr_read_data2[2]
port 155 nsew signal input
rlabel metal2 s 191010 199200 191066 200000 6 instr_read_data2[30]
port 156 nsew signal input
rlabel metal2 s 193954 199200 194010 200000 6 instr_read_data2[31]
port 157 nsew signal input
rlabel metal2 s 103058 199200 103114 200000 6 instr_read_data2[3]
port 158 nsew signal input
rlabel metal2 s 107474 199200 107530 200000 6 instr_read_data2[4]
port 159 nsew signal input
rlabel metal2 s 111522 199200 111578 200000 6 instr_read_data2[5]
port 160 nsew signal input
rlabel metal2 s 115570 199200 115626 200000 6 instr_read_data2[6]
port 161 nsew signal input
rlabel metal2 s 119618 199200 119674 200000 6 instr_read_data2[7]
port 162 nsew signal input
rlabel metal2 s 123298 199200 123354 200000 6 instr_read_data2[8]
port 163 nsew signal input
rlabel metal2 s 126610 199200 126666 200000 6 instr_read_data2[9]
port 164 nsew signal input
rlabel metal2 s 90178 199200 90234 200000 6 instr_read_data3[0]
port 165 nsew signal input
rlabel metal2 s 130290 199200 130346 200000 6 instr_read_data3[10]
port 166 nsew signal input
rlabel metal2 s 133602 199200 133658 200000 6 instr_read_data3[11]
port 167 nsew signal input
rlabel metal2 s 136914 199200 136970 200000 6 instr_read_data3[12]
port 168 nsew signal input
rlabel metal2 s 140226 199200 140282 200000 6 instr_read_data3[13]
port 169 nsew signal input
rlabel metal2 s 143538 199200 143594 200000 6 instr_read_data3[14]
port 170 nsew signal input
rlabel metal2 s 146850 199200 146906 200000 6 instr_read_data3[15]
port 171 nsew signal input
rlabel metal2 s 150162 199200 150218 200000 6 instr_read_data3[16]
port 172 nsew signal input
rlabel metal2 s 153106 199200 153162 200000 6 instr_read_data3[17]
port 173 nsew signal input
rlabel metal2 s 156050 199200 156106 200000 6 instr_read_data3[18]
port 174 nsew signal input
rlabel metal2 s 158994 199200 159050 200000 6 instr_read_data3[19]
port 175 nsew signal input
rlabel metal2 s 94594 199200 94650 200000 6 instr_read_data3[1]
port 176 nsew signal input
rlabel metal2 s 161938 199200 161994 200000 6 instr_read_data3[20]
port 177 nsew signal input
rlabel metal2 s 164882 199200 164938 200000 6 instr_read_data3[21]
port 178 nsew signal input
rlabel metal2 s 167826 199200 167882 200000 6 instr_read_data3[22]
port 179 nsew signal input
rlabel metal2 s 170770 199200 170826 200000 6 instr_read_data3[23]
port 180 nsew signal input
rlabel metal2 s 173714 199200 173770 200000 6 instr_read_data3[24]
port 181 nsew signal input
rlabel metal2 s 176658 199200 176714 200000 6 instr_read_data3[25]
port 182 nsew signal input
rlabel metal2 s 179602 199200 179658 200000 6 instr_read_data3[26]
port 183 nsew signal input
rlabel metal2 s 182546 199200 182602 200000 6 instr_read_data3[27]
port 184 nsew signal input
rlabel metal2 s 185490 199200 185546 200000 6 instr_read_data3[28]
port 185 nsew signal input
rlabel metal2 s 188434 199200 188490 200000 6 instr_read_data3[29]
port 186 nsew signal input
rlabel metal2 s 99010 199200 99066 200000 6 instr_read_data3[2]
port 187 nsew signal input
rlabel metal2 s 191378 199200 191434 200000 6 instr_read_data3[30]
port 188 nsew signal input
rlabel metal2 s 194322 199200 194378 200000 6 instr_read_data3[31]
port 189 nsew signal input
rlabel metal2 s 103426 199200 103482 200000 6 instr_read_data3[3]
port 190 nsew signal input
rlabel metal2 s 107842 199200 107898 200000 6 instr_read_data3[4]
port 191 nsew signal input
rlabel metal2 s 111890 199200 111946 200000 6 instr_read_data3[5]
port 192 nsew signal input
rlabel metal2 s 115938 199200 115994 200000 6 instr_read_data3[6]
port 193 nsew signal input
rlabel metal2 s 119986 199200 120042 200000 6 instr_read_data3[7]
port 194 nsew signal input
rlabel metal2 s 123666 199200 123722 200000 6 instr_read_data3[8]
port 195 nsew signal input
rlabel metal2 s 126978 199200 127034 200000 6 instr_read_data3[9]
port 196 nsew signal input
rlabel metal2 s 90546 199200 90602 200000 6 instr_read_data4[0]
port 197 nsew signal input
rlabel metal2 s 130658 199200 130714 200000 6 instr_read_data4[10]
port 198 nsew signal input
rlabel metal2 s 133970 199200 134026 200000 6 instr_read_data4[11]
port 199 nsew signal input
rlabel metal2 s 137282 199200 137338 200000 6 instr_read_data4[12]
port 200 nsew signal input
rlabel metal2 s 140594 199200 140650 200000 6 instr_read_data4[13]
port 201 nsew signal input
rlabel metal2 s 143906 199200 143962 200000 6 instr_read_data4[14]
port 202 nsew signal input
rlabel metal2 s 147218 199200 147274 200000 6 instr_read_data4[15]
port 203 nsew signal input
rlabel metal2 s 150530 199200 150586 200000 6 instr_read_data4[16]
port 204 nsew signal input
rlabel metal2 s 153474 199200 153530 200000 6 instr_read_data4[17]
port 205 nsew signal input
rlabel metal2 s 156418 199200 156474 200000 6 instr_read_data4[18]
port 206 nsew signal input
rlabel metal2 s 159362 199200 159418 200000 6 instr_read_data4[19]
port 207 nsew signal input
rlabel metal2 s 94962 199200 95018 200000 6 instr_read_data4[1]
port 208 nsew signal input
rlabel metal2 s 162306 199200 162362 200000 6 instr_read_data4[20]
port 209 nsew signal input
rlabel metal2 s 165250 199200 165306 200000 6 instr_read_data4[21]
port 210 nsew signal input
rlabel metal2 s 168194 199200 168250 200000 6 instr_read_data4[22]
port 211 nsew signal input
rlabel metal2 s 171138 199200 171194 200000 6 instr_read_data4[23]
port 212 nsew signal input
rlabel metal2 s 174082 199200 174138 200000 6 instr_read_data4[24]
port 213 nsew signal input
rlabel metal2 s 177026 199200 177082 200000 6 instr_read_data4[25]
port 214 nsew signal input
rlabel metal2 s 179970 199200 180026 200000 6 instr_read_data4[26]
port 215 nsew signal input
rlabel metal2 s 182914 199200 182970 200000 6 instr_read_data4[27]
port 216 nsew signal input
rlabel metal2 s 185858 199200 185914 200000 6 instr_read_data4[28]
port 217 nsew signal input
rlabel metal2 s 188802 199200 188858 200000 6 instr_read_data4[29]
port 218 nsew signal input
rlabel metal2 s 99378 199200 99434 200000 6 instr_read_data4[2]
port 219 nsew signal input
rlabel metal2 s 191746 199200 191802 200000 6 instr_read_data4[30]
port 220 nsew signal input
rlabel metal2 s 194690 199200 194746 200000 6 instr_read_data4[31]
port 221 nsew signal input
rlabel metal2 s 103794 199200 103850 200000 6 instr_read_data4[3]
port 222 nsew signal input
rlabel metal2 s 108210 199200 108266 200000 6 instr_read_data4[4]
port 223 nsew signal input
rlabel metal2 s 112258 199200 112314 200000 6 instr_read_data4[5]
port 224 nsew signal input
rlabel metal2 s 116306 199200 116362 200000 6 instr_read_data4[6]
port 225 nsew signal input
rlabel metal2 s 120354 199200 120410 200000 6 instr_read_data4[7]
port 226 nsew signal input
rlabel metal2 s 124034 199200 124090 200000 6 instr_read_data4[8]
port 227 nsew signal input
rlabel metal2 s 127346 199200 127402 200000 6 instr_read_data4[9]
port 228 nsew signal input
rlabel metal2 s 90914 199200 90970 200000 6 instr_read_data5[0]
port 229 nsew signal input
rlabel metal2 s 131026 199200 131082 200000 6 instr_read_data5[10]
port 230 nsew signal input
rlabel metal2 s 134338 199200 134394 200000 6 instr_read_data5[11]
port 231 nsew signal input
rlabel metal2 s 137650 199200 137706 200000 6 instr_read_data5[12]
port 232 nsew signal input
rlabel metal2 s 140962 199200 141018 200000 6 instr_read_data5[13]
port 233 nsew signal input
rlabel metal2 s 144274 199200 144330 200000 6 instr_read_data5[14]
port 234 nsew signal input
rlabel metal2 s 147586 199200 147642 200000 6 instr_read_data5[15]
port 235 nsew signal input
rlabel metal2 s 150898 199200 150954 200000 6 instr_read_data5[16]
port 236 nsew signal input
rlabel metal2 s 153842 199200 153898 200000 6 instr_read_data5[17]
port 237 nsew signal input
rlabel metal2 s 156786 199200 156842 200000 6 instr_read_data5[18]
port 238 nsew signal input
rlabel metal2 s 159730 199200 159786 200000 6 instr_read_data5[19]
port 239 nsew signal input
rlabel metal2 s 95330 199200 95386 200000 6 instr_read_data5[1]
port 240 nsew signal input
rlabel metal2 s 162674 199200 162730 200000 6 instr_read_data5[20]
port 241 nsew signal input
rlabel metal2 s 165618 199200 165674 200000 6 instr_read_data5[21]
port 242 nsew signal input
rlabel metal2 s 168562 199200 168618 200000 6 instr_read_data5[22]
port 243 nsew signal input
rlabel metal2 s 171506 199200 171562 200000 6 instr_read_data5[23]
port 244 nsew signal input
rlabel metal2 s 174450 199200 174506 200000 6 instr_read_data5[24]
port 245 nsew signal input
rlabel metal2 s 177394 199200 177450 200000 6 instr_read_data5[25]
port 246 nsew signal input
rlabel metal2 s 180338 199200 180394 200000 6 instr_read_data5[26]
port 247 nsew signal input
rlabel metal2 s 183282 199200 183338 200000 6 instr_read_data5[27]
port 248 nsew signal input
rlabel metal2 s 186226 199200 186282 200000 6 instr_read_data5[28]
port 249 nsew signal input
rlabel metal2 s 189170 199200 189226 200000 6 instr_read_data5[29]
port 250 nsew signal input
rlabel metal2 s 99746 199200 99802 200000 6 instr_read_data5[2]
port 251 nsew signal input
rlabel metal2 s 192114 199200 192170 200000 6 instr_read_data5[30]
port 252 nsew signal input
rlabel metal2 s 195058 199200 195114 200000 6 instr_read_data5[31]
port 253 nsew signal input
rlabel metal2 s 104162 199200 104218 200000 6 instr_read_data5[3]
port 254 nsew signal input
rlabel metal2 s 108578 199200 108634 200000 6 instr_read_data5[4]
port 255 nsew signal input
rlabel metal2 s 112626 199200 112682 200000 6 instr_read_data5[5]
port 256 nsew signal input
rlabel metal2 s 116674 199200 116730 200000 6 instr_read_data5[6]
port 257 nsew signal input
rlabel metal2 s 120722 199200 120778 200000 6 instr_read_data5[7]
port 258 nsew signal input
rlabel metal2 s 124402 199200 124458 200000 6 instr_read_data5[8]
port 259 nsew signal input
rlabel metal2 s 127714 199200 127770 200000 6 instr_read_data5[9]
port 260 nsew signal input
rlabel metal2 s 91282 199200 91338 200000 6 instr_read_data6[0]
port 261 nsew signal input
rlabel metal2 s 131394 199200 131450 200000 6 instr_read_data6[10]
port 262 nsew signal input
rlabel metal2 s 134706 199200 134762 200000 6 instr_read_data6[11]
port 263 nsew signal input
rlabel metal2 s 138018 199200 138074 200000 6 instr_read_data6[12]
port 264 nsew signal input
rlabel metal2 s 141330 199200 141386 200000 6 instr_read_data6[13]
port 265 nsew signal input
rlabel metal2 s 144642 199200 144698 200000 6 instr_read_data6[14]
port 266 nsew signal input
rlabel metal2 s 147954 199200 148010 200000 6 instr_read_data6[15]
port 267 nsew signal input
rlabel metal2 s 151266 199200 151322 200000 6 instr_read_data6[16]
port 268 nsew signal input
rlabel metal2 s 154210 199200 154266 200000 6 instr_read_data6[17]
port 269 nsew signal input
rlabel metal2 s 157154 199200 157210 200000 6 instr_read_data6[18]
port 270 nsew signal input
rlabel metal2 s 160098 199200 160154 200000 6 instr_read_data6[19]
port 271 nsew signal input
rlabel metal2 s 95698 199200 95754 200000 6 instr_read_data6[1]
port 272 nsew signal input
rlabel metal2 s 163042 199200 163098 200000 6 instr_read_data6[20]
port 273 nsew signal input
rlabel metal2 s 165986 199200 166042 200000 6 instr_read_data6[21]
port 274 nsew signal input
rlabel metal2 s 168930 199200 168986 200000 6 instr_read_data6[22]
port 275 nsew signal input
rlabel metal2 s 171874 199200 171930 200000 6 instr_read_data6[23]
port 276 nsew signal input
rlabel metal2 s 174818 199200 174874 200000 6 instr_read_data6[24]
port 277 nsew signal input
rlabel metal2 s 177762 199200 177818 200000 6 instr_read_data6[25]
port 278 nsew signal input
rlabel metal2 s 180706 199200 180762 200000 6 instr_read_data6[26]
port 279 nsew signal input
rlabel metal2 s 183650 199200 183706 200000 6 instr_read_data6[27]
port 280 nsew signal input
rlabel metal2 s 186594 199200 186650 200000 6 instr_read_data6[28]
port 281 nsew signal input
rlabel metal2 s 189538 199200 189594 200000 6 instr_read_data6[29]
port 282 nsew signal input
rlabel metal2 s 100114 199200 100170 200000 6 instr_read_data6[2]
port 283 nsew signal input
rlabel metal2 s 192482 199200 192538 200000 6 instr_read_data6[30]
port 284 nsew signal input
rlabel metal2 s 195426 199200 195482 200000 6 instr_read_data6[31]
port 285 nsew signal input
rlabel metal2 s 104530 199200 104586 200000 6 instr_read_data6[3]
port 286 nsew signal input
rlabel metal2 s 108946 199200 109002 200000 6 instr_read_data6[4]
port 287 nsew signal input
rlabel metal2 s 112994 199200 113050 200000 6 instr_read_data6[5]
port 288 nsew signal input
rlabel metal2 s 117042 199200 117098 200000 6 instr_read_data6[6]
port 289 nsew signal input
rlabel metal2 s 121090 199200 121146 200000 6 instr_read_data6[7]
port 290 nsew signal input
rlabel metal2 s 124770 199200 124826 200000 6 instr_read_data6[8]
port 291 nsew signal input
rlabel metal2 s 128082 199200 128138 200000 6 instr_read_data6[9]
port 292 nsew signal input
rlabel metal2 s 91650 199200 91706 200000 6 instr_read_data7[0]
port 293 nsew signal input
rlabel metal2 s 131762 199200 131818 200000 6 instr_read_data7[10]
port 294 nsew signal input
rlabel metal2 s 135074 199200 135130 200000 6 instr_read_data7[11]
port 295 nsew signal input
rlabel metal2 s 138386 199200 138442 200000 6 instr_read_data7[12]
port 296 nsew signal input
rlabel metal2 s 141698 199200 141754 200000 6 instr_read_data7[13]
port 297 nsew signal input
rlabel metal2 s 145010 199200 145066 200000 6 instr_read_data7[14]
port 298 nsew signal input
rlabel metal2 s 148322 199200 148378 200000 6 instr_read_data7[15]
port 299 nsew signal input
rlabel metal2 s 151634 199200 151690 200000 6 instr_read_data7[16]
port 300 nsew signal input
rlabel metal2 s 154578 199200 154634 200000 6 instr_read_data7[17]
port 301 nsew signal input
rlabel metal2 s 157522 199200 157578 200000 6 instr_read_data7[18]
port 302 nsew signal input
rlabel metal2 s 160466 199200 160522 200000 6 instr_read_data7[19]
port 303 nsew signal input
rlabel metal2 s 96066 199200 96122 200000 6 instr_read_data7[1]
port 304 nsew signal input
rlabel metal2 s 163410 199200 163466 200000 6 instr_read_data7[20]
port 305 nsew signal input
rlabel metal2 s 166354 199200 166410 200000 6 instr_read_data7[21]
port 306 nsew signal input
rlabel metal2 s 169298 199200 169354 200000 6 instr_read_data7[22]
port 307 nsew signal input
rlabel metal2 s 172242 199200 172298 200000 6 instr_read_data7[23]
port 308 nsew signal input
rlabel metal2 s 175186 199200 175242 200000 6 instr_read_data7[24]
port 309 nsew signal input
rlabel metal2 s 178130 199200 178186 200000 6 instr_read_data7[25]
port 310 nsew signal input
rlabel metal2 s 181074 199200 181130 200000 6 instr_read_data7[26]
port 311 nsew signal input
rlabel metal2 s 184018 199200 184074 200000 6 instr_read_data7[27]
port 312 nsew signal input
rlabel metal2 s 186962 199200 187018 200000 6 instr_read_data7[28]
port 313 nsew signal input
rlabel metal2 s 189906 199200 189962 200000 6 instr_read_data7[29]
port 314 nsew signal input
rlabel metal2 s 100482 199200 100538 200000 6 instr_read_data7[2]
port 315 nsew signal input
rlabel metal2 s 192850 199200 192906 200000 6 instr_read_data7[30]
port 316 nsew signal input
rlabel metal2 s 195794 199200 195850 200000 6 instr_read_data7[31]
port 317 nsew signal input
rlabel metal2 s 104898 199200 104954 200000 6 instr_read_data7[3]
port 318 nsew signal input
rlabel metal2 s 109314 199200 109370 200000 6 instr_read_data7[4]
port 319 nsew signal input
rlabel metal2 s 113362 199200 113418 200000 6 instr_read_data7[5]
port 320 nsew signal input
rlabel metal2 s 117410 199200 117466 200000 6 instr_read_data7[6]
port 321 nsew signal input
rlabel metal2 s 121458 199200 121514 200000 6 instr_read_data7[7]
port 322 nsew signal input
rlabel metal2 s 125138 199200 125194 200000 6 instr_read_data7[8]
port 323 nsew signal input
rlabel metal2 s 128450 199200 128506 200000 6 instr_read_data7[9]
port 324 nsew signal input
rlabel metal2 s 92018 199200 92074 200000 6 instr_wmask[0]
port 325 nsew signal output
rlabel metal2 s 96434 199200 96490 200000 6 instr_wmask[1]
port 326 nsew signal output
rlabel metal2 s 100850 199200 100906 200000 6 instr_wmask[2]
port 327 nsew signal output
rlabel metal2 s 105266 199200 105322 200000 6 instr_wmask[3]
port 328 nsew signal output
rlabel metal2 s 92386 199200 92442 200000 6 instr_write_data[0]
port 329 nsew signal output
rlabel metal2 s 132130 199200 132186 200000 6 instr_write_data[10]
port 330 nsew signal output
rlabel metal2 s 135442 199200 135498 200000 6 instr_write_data[11]
port 331 nsew signal output
rlabel metal2 s 138754 199200 138810 200000 6 instr_write_data[12]
port 332 nsew signal output
rlabel metal2 s 142066 199200 142122 200000 6 instr_write_data[13]
port 333 nsew signal output
rlabel metal2 s 145378 199200 145434 200000 6 instr_write_data[14]
port 334 nsew signal output
rlabel metal2 s 148690 199200 148746 200000 6 instr_write_data[15]
port 335 nsew signal output
rlabel metal2 s 96802 199200 96858 200000 6 instr_write_data[1]
port 336 nsew signal output
rlabel metal2 s 101218 199200 101274 200000 6 instr_write_data[2]
port 337 nsew signal output
rlabel metal2 s 105634 199200 105690 200000 6 instr_write_data[3]
port 338 nsew signal output
rlabel metal2 s 109682 199200 109738 200000 6 instr_write_data[4]
port 339 nsew signal output
rlabel metal2 s 113730 199200 113786 200000 6 instr_write_data[5]
port 340 nsew signal output
rlabel metal2 s 117778 199200 117834 200000 6 instr_write_data[6]
port 341 nsew signal output
rlabel metal2 s 121826 199200 121882 200000 6 instr_write_data[7]
port 342 nsew signal output
rlabel metal2 s 125506 199200 125562 200000 6 instr_write_data[8]
port 343 nsew signal output
rlabel metal2 s 128818 199200 128874 200000 6 instr_write_data[9]
port 344 nsew signal output
rlabel metal2 s 196162 199200 196218 200000 6 instrw_enb
port 345 nsew signal output
rlabel metal2 s 3698 199200 3754 200000 6 io_in[0]
port 346 nsew signal input
rlabel metal2 s 14738 199200 14794 200000 6 io_in[10]
port 347 nsew signal input
rlabel metal2 s 15842 199200 15898 200000 6 io_in[11]
port 348 nsew signal input
rlabel metal2 s 16946 199200 17002 200000 6 io_in[12]
port 349 nsew signal input
rlabel metal2 s 18050 199200 18106 200000 6 io_in[13]
port 350 nsew signal input
rlabel metal2 s 19154 199200 19210 200000 6 io_in[14]
port 351 nsew signal input
rlabel metal2 s 20258 199200 20314 200000 6 io_in[15]
port 352 nsew signal input
rlabel metal2 s 21362 199200 21418 200000 6 io_in[16]
port 353 nsew signal input
rlabel metal2 s 22466 199200 22522 200000 6 io_in[17]
port 354 nsew signal input
rlabel metal2 s 23570 199200 23626 200000 6 io_in[18]
port 355 nsew signal input
rlabel metal2 s 24674 199200 24730 200000 6 io_in[19]
port 356 nsew signal input
rlabel metal2 s 4802 199200 4858 200000 6 io_in[1]
port 357 nsew signal input
rlabel metal2 s 25778 199200 25834 200000 6 io_in[20]
port 358 nsew signal input
rlabel metal2 s 26882 199200 26938 200000 6 io_in[21]
port 359 nsew signal input
rlabel metal2 s 27986 199200 28042 200000 6 io_in[22]
port 360 nsew signal input
rlabel metal2 s 29090 199200 29146 200000 6 io_in[23]
port 361 nsew signal input
rlabel metal2 s 30194 199200 30250 200000 6 io_in[24]
port 362 nsew signal input
rlabel metal2 s 31298 199200 31354 200000 6 io_in[25]
port 363 nsew signal input
rlabel metal2 s 32402 199200 32458 200000 6 io_in[26]
port 364 nsew signal input
rlabel metal2 s 33506 199200 33562 200000 6 io_in[27]
port 365 nsew signal input
rlabel metal2 s 34610 199200 34666 200000 6 io_in[28]
port 366 nsew signal input
rlabel metal2 s 35714 199200 35770 200000 6 io_in[29]
port 367 nsew signal input
rlabel metal2 s 5906 199200 5962 200000 6 io_in[2]
port 368 nsew signal input
rlabel metal2 s 36818 199200 36874 200000 6 io_in[30]
port 369 nsew signal input
rlabel metal2 s 37922 199200 37978 200000 6 io_in[31]
port 370 nsew signal input
rlabel metal2 s 39026 199200 39082 200000 6 io_in[32]
port 371 nsew signal input
rlabel metal2 s 40130 199200 40186 200000 6 io_in[33]
port 372 nsew signal input
rlabel metal2 s 41234 199200 41290 200000 6 io_in[34]
port 373 nsew signal input
rlabel metal2 s 42338 199200 42394 200000 6 io_in[35]
port 374 nsew signal input
rlabel metal2 s 43442 199200 43498 200000 6 io_in[36]
port 375 nsew signal input
rlabel metal2 s 44546 199200 44602 200000 6 io_in[37]
port 376 nsew signal input
rlabel metal2 s 7010 199200 7066 200000 6 io_in[3]
port 377 nsew signal input
rlabel metal2 s 8114 199200 8170 200000 6 io_in[4]
port 378 nsew signal input
rlabel metal2 s 9218 199200 9274 200000 6 io_in[5]
port 379 nsew signal input
rlabel metal2 s 10322 199200 10378 200000 6 io_in[6]
port 380 nsew signal input
rlabel metal2 s 11426 199200 11482 200000 6 io_in[7]
port 381 nsew signal input
rlabel metal2 s 12530 199200 12586 200000 6 io_in[8]
port 382 nsew signal input
rlabel metal2 s 13634 199200 13690 200000 6 io_in[9]
port 383 nsew signal input
rlabel metal2 s 4066 199200 4122 200000 6 io_oeb[0]
port 384 nsew signal output
rlabel metal2 s 15106 199200 15162 200000 6 io_oeb[10]
port 385 nsew signal output
rlabel metal2 s 16210 199200 16266 200000 6 io_oeb[11]
port 386 nsew signal output
rlabel metal2 s 17314 199200 17370 200000 6 io_oeb[12]
port 387 nsew signal output
rlabel metal2 s 18418 199200 18474 200000 6 io_oeb[13]
port 388 nsew signal output
rlabel metal2 s 19522 199200 19578 200000 6 io_oeb[14]
port 389 nsew signal output
rlabel metal2 s 20626 199200 20682 200000 6 io_oeb[15]
port 390 nsew signal output
rlabel metal2 s 21730 199200 21786 200000 6 io_oeb[16]
port 391 nsew signal output
rlabel metal2 s 22834 199200 22890 200000 6 io_oeb[17]
port 392 nsew signal output
rlabel metal2 s 23938 199200 23994 200000 6 io_oeb[18]
port 393 nsew signal output
rlabel metal2 s 25042 199200 25098 200000 6 io_oeb[19]
port 394 nsew signal output
rlabel metal2 s 5170 199200 5226 200000 6 io_oeb[1]
port 395 nsew signal output
rlabel metal2 s 26146 199200 26202 200000 6 io_oeb[20]
port 396 nsew signal output
rlabel metal2 s 27250 199200 27306 200000 6 io_oeb[21]
port 397 nsew signal output
rlabel metal2 s 28354 199200 28410 200000 6 io_oeb[22]
port 398 nsew signal output
rlabel metal2 s 29458 199200 29514 200000 6 io_oeb[23]
port 399 nsew signal output
rlabel metal2 s 30562 199200 30618 200000 6 io_oeb[24]
port 400 nsew signal output
rlabel metal2 s 31666 199200 31722 200000 6 io_oeb[25]
port 401 nsew signal output
rlabel metal2 s 32770 199200 32826 200000 6 io_oeb[26]
port 402 nsew signal output
rlabel metal2 s 33874 199200 33930 200000 6 io_oeb[27]
port 403 nsew signal output
rlabel metal2 s 34978 199200 35034 200000 6 io_oeb[28]
port 404 nsew signal output
rlabel metal2 s 36082 199200 36138 200000 6 io_oeb[29]
port 405 nsew signal output
rlabel metal2 s 6274 199200 6330 200000 6 io_oeb[2]
port 406 nsew signal output
rlabel metal2 s 37186 199200 37242 200000 6 io_oeb[30]
port 407 nsew signal output
rlabel metal2 s 38290 199200 38346 200000 6 io_oeb[31]
port 408 nsew signal output
rlabel metal2 s 39394 199200 39450 200000 6 io_oeb[32]
port 409 nsew signal output
rlabel metal2 s 40498 199200 40554 200000 6 io_oeb[33]
port 410 nsew signal output
rlabel metal2 s 41602 199200 41658 200000 6 io_oeb[34]
port 411 nsew signal output
rlabel metal2 s 42706 199200 42762 200000 6 io_oeb[35]
port 412 nsew signal output
rlabel metal2 s 43810 199200 43866 200000 6 io_oeb[36]
port 413 nsew signal output
rlabel metal2 s 44914 199200 44970 200000 6 io_oeb[37]
port 414 nsew signal output
rlabel metal2 s 7378 199200 7434 200000 6 io_oeb[3]
port 415 nsew signal output
rlabel metal2 s 8482 199200 8538 200000 6 io_oeb[4]
port 416 nsew signal output
rlabel metal2 s 9586 199200 9642 200000 6 io_oeb[5]
port 417 nsew signal output
rlabel metal2 s 10690 199200 10746 200000 6 io_oeb[6]
port 418 nsew signal output
rlabel metal2 s 11794 199200 11850 200000 6 io_oeb[7]
port 419 nsew signal output
rlabel metal2 s 12898 199200 12954 200000 6 io_oeb[8]
port 420 nsew signal output
rlabel metal2 s 14002 199200 14058 200000 6 io_oeb[9]
port 421 nsew signal output
rlabel metal2 s 4434 199200 4490 200000 6 io_out[0]
port 422 nsew signal output
rlabel metal2 s 15474 199200 15530 200000 6 io_out[10]
port 423 nsew signal output
rlabel metal2 s 16578 199200 16634 200000 6 io_out[11]
port 424 nsew signal output
rlabel metal2 s 17682 199200 17738 200000 6 io_out[12]
port 425 nsew signal output
rlabel metal2 s 18786 199200 18842 200000 6 io_out[13]
port 426 nsew signal output
rlabel metal2 s 19890 199200 19946 200000 6 io_out[14]
port 427 nsew signal output
rlabel metal2 s 20994 199200 21050 200000 6 io_out[15]
port 428 nsew signal output
rlabel metal2 s 22098 199200 22154 200000 6 io_out[16]
port 429 nsew signal output
rlabel metal2 s 23202 199200 23258 200000 6 io_out[17]
port 430 nsew signal output
rlabel metal2 s 24306 199200 24362 200000 6 io_out[18]
port 431 nsew signal output
rlabel metal2 s 25410 199200 25466 200000 6 io_out[19]
port 432 nsew signal output
rlabel metal2 s 5538 199200 5594 200000 6 io_out[1]
port 433 nsew signal output
rlabel metal2 s 26514 199200 26570 200000 6 io_out[20]
port 434 nsew signal output
rlabel metal2 s 27618 199200 27674 200000 6 io_out[21]
port 435 nsew signal output
rlabel metal2 s 28722 199200 28778 200000 6 io_out[22]
port 436 nsew signal output
rlabel metal2 s 29826 199200 29882 200000 6 io_out[23]
port 437 nsew signal output
rlabel metal2 s 30930 199200 30986 200000 6 io_out[24]
port 438 nsew signal output
rlabel metal2 s 32034 199200 32090 200000 6 io_out[25]
port 439 nsew signal output
rlabel metal2 s 33138 199200 33194 200000 6 io_out[26]
port 440 nsew signal output
rlabel metal2 s 34242 199200 34298 200000 6 io_out[27]
port 441 nsew signal output
rlabel metal2 s 35346 199200 35402 200000 6 io_out[28]
port 442 nsew signal output
rlabel metal2 s 36450 199200 36506 200000 6 io_out[29]
port 443 nsew signal output
rlabel metal2 s 6642 199200 6698 200000 6 io_out[2]
port 444 nsew signal output
rlabel metal2 s 37554 199200 37610 200000 6 io_out[30]
port 445 nsew signal output
rlabel metal2 s 38658 199200 38714 200000 6 io_out[31]
port 446 nsew signal output
rlabel metal2 s 39762 199200 39818 200000 6 io_out[32]
port 447 nsew signal output
rlabel metal2 s 40866 199200 40922 200000 6 io_out[33]
port 448 nsew signal output
rlabel metal2 s 41970 199200 42026 200000 6 io_out[34]
port 449 nsew signal output
rlabel metal2 s 43074 199200 43130 200000 6 io_out[35]
port 450 nsew signal output
rlabel metal2 s 44178 199200 44234 200000 6 io_out[36]
port 451 nsew signal output
rlabel metal2 s 45282 199200 45338 200000 6 io_out[37]
port 452 nsew signal output
rlabel metal2 s 7746 199200 7802 200000 6 io_out[3]
port 453 nsew signal output
rlabel metal2 s 8850 199200 8906 200000 6 io_out[4]
port 454 nsew signal output
rlabel metal2 s 9954 199200 10010 200000 6 io_out[5]
port 455 nsew signal output
rlabel metal2 s 11058 199200 11114 200000 6 io_out[6]
port 456 nsew signal output
rlabel metal2 s 12162 199200 12218 200000 6 io_out[7]
port 457 nsew signal output
rlabel metal2 s 13266 199200 13322 200000 6 io_out[8]
port 458 nsew signal output
rlabel metal2 s 14370 199200 14426 200000 6 io_out[9]
port 459 nsew signal output
rlabel metal2 s 184110 0 184166 800 6 irq[0]
port 460 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 irq[1]
port 461 nsew signal output
rlabel metal2 s 186870 0 186926 800 6 irq[2]
port 462 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 la_data_in
port 463 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 la_data_out[0]
port 464 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[100]
port 465 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[101]
port 466 nsew signal output
rlabel metal2 s 148230 0 148286 800 6 la_data_out[102]
port 467 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[103]
port 468 nsew signal output
rlabel metal2 s 150990 0 151046 800 6 la_data_out[104]
port 469 nsew signal output
rlabel metal2 s 152370 0 152426 800 6 la_data_out[105]
port 470 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[106]
port 471 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[107]
port 472 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[108]
port 473 nsew signal output
rlabel metal2 s 157890 0 157946 800 6 la_data_out[109]
port 474 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 la_data_out[10]
port 475 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 la_data_out[110]
port 476 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[111]
port 477 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[112]
port 478 nsew signal output
rlabel metal2 s 163410 0 163466 800 6 la_data_out[113]
port 479 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 la_data_out[114]
port 480 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 la_data_out[115]
port 481 nsew signal output
rlabel metal2 s 167550 0 167606 800 6 la_data_out[116]
port 482 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[117]
port 483 nsew signal output
rlabel metal2 s 170310 0 170366 800 6 la_data_out[118]
port 484 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 la_data_out[119]
port 485 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 la_data_out[11]
port 486 nsew signal output
rlabel metal2 s 173070 0 173126 800 6 la_data_out[120]
port 487 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 la_data_out[121]
port 488 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[122]
port 489 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[123]
port 490 nsew signal output
rlabel metal2 s 178590 0 178646 800 6 la_data_out[124]
port 491 nsew signal output
rlabel metal2 s 179970 0 180026 800 6 la_data_out[125]
port 492 nsew signal output
rlabel metal2 s 181350 0 181406 800 6 la_data_out[126]
port 493 nsew signal output
rlabel metal2 s 182730 0 182786 800 6 la_data_out[127]
port 494 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 la_data_out[12]
port 495 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 la_data_out[13]
port 496 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 la_data_out[14]
port 497 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 la_data_out[15]
port 498 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_out[16]
port 499 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 la_data_out[17]
port 500 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 la_data_out[18]
port 501 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 la_data_out[19]
port 502 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 la_data_out[1]
port 503 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_data_out[20]
port 504 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 la_data_out[21]
port 505 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 la_data_out[22]
port 506 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 la_data_out[23]
port 507 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[24]
port 508 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[25]
port 509 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 la_data_out[26]
port 510 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[27]
port 511 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[28]
port 512 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[29]
port 513 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 la_data_out[2]
port 514 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[30]
port 515 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 la_data_out[31]
port 516 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[32]
port 517 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 la_data_out[33]
port 518 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 la_data_out[34]
port 519 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[35]
port 520 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[36]
port 521 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[37]
port 522 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 la_data_out[38]
port 523 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[39]
port 524 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 la_data_out[3]
port 525 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 la_data_out[40]
port 526 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[41]
port 527 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[42]
port 528 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[43]
port 529 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[44]
port 530 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[45]
port 531 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 la_data_out[46]
port 532 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[47]
port 533 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[48]
port 534 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 la_data_out[49]
port 535 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 la_data_out[4]
port 536 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[50]
port 537 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[51]
port 538 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[52]
port 539 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[53]
port 540 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[54]
port 541 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[55]
port 542 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[56]
port 543 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[57]
port 544 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[58]
port 545 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[59]
port 546 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 la_data_out[5]
port 547 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[60]
port 548 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[61]
port 549 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[62]
port 550 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[63]
port 551 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[64]
port 552 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[65]
port 553 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[66]
port 554 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[67]
port 555 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[68]
port 556 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 la_data_out[69]
port 557 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 la_data_out[6]
port 558 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 la_data_out[70]
port 559 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 la_data_out[71]
port 560 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[72]
port 561 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[73]
port 562 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 la_data_out[74]
port 563 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[75]
port 564 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 la_data_out[76]
port 565 nsew signal output
rlabel metal2 s 113730 0 113786 800 6 la_data_out[77]
port 566 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[78]
port 567 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[79]
port 568 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 la_data_out[7]
port 569 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[80]
port 570 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 la_data_out[81]
port 571 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 la_data_out[82]
port 572 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[83]
port 573 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[84]
port 574 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 la_data_out[85]
port 575 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[86]
port 576 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[87]
port 577 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[88]
port 578 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[89]
port 579 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 la_data_out[8]
port 580 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 la_data_out[90]
port 581 nsew signal output
rlabel metal2 s 133050 0 133106 800 6 la_data_out[91]
port 582 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[92]
port 583 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[93]
port 584 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[94]
port 585 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[95]
port 586 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[96]
port 587 nsew signal output
rlabel metal2 s 141330 0 141386 800 6 la_data_out[97]
port 588 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 la_data_out[98]
port 589 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 la_data_out[99]
port 590 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 la_data_out[9]
port 591 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 la_oenb
port 592 nsew signal input
rlabel metal2 s 197910 0 197966 800 6 low
port 593 nsew signal output
rlabel metal2 s 189630 0 189686 800 6 reset
port 594 nsew signal output
rlabel metal2 s 191010 0 191066 800 6 start
port 595 nsew signal output
rlabel metal2 s 46018 199200 46074 200000 6 uP_data_mem_addr[0]
port 596 nsew signal input
rlabel metal2 s 47858 199200 47914 200000 6 uP_data_mem_addr[1]
port 597 nsew signal input
rlabel metal2 s 49698 199200 49754 200000 6 uP_data_mem_addr[2]
port 598 nsew signal input
rlabel metal2 s 51538 199200 51594 200000 6 uP_data_mem_addr[3]
port 599 nsew signal input
rlabel metal2 s 53378 199200 53434 200000 6 uP_data_mem_addr[4]
port 600 nsew signal input
rlabel metal2 s 55218 199200 55274 200000 6 uP_data_mem_addr[5]
port 601 nsew signal input
rlabel metal2 s 57058 199200 57114 200000 6 uP_data_mem_addr[6]
port 602 nsew signal input
rlabel metal2 s 58898 199200 58954 200000 6 uP_data_mem_addr[7]
port 603 nsew signal input
rlabel metal2 s 45650 199200 45706 200000 6 uP_dataw_en
port 604 nsew signal input
rlabel metal2 s 46386 199200 46442 200000 6 uP_instr[0]
port 605 nsew signal output
rlabel metal2 s 63682 199200 63738 200000 6 uP_instr[10]
port 606 nsew signal output
rlabel metal2 s 65154 199200 65210 200000 6 uP_instr[11]
port 607 nsew signal output
rlabel metal2 s 66626 199200 66682 200000 6 uP_instr[12]
port 608 nsew signal output
rlabel metal2 s 68098 199200 68154 200000 6 uP_instr[13]
port 609 nsew signal output
rlabel metal2 s 69202 199200 69258 200000 6 uP_instr[14]
port 610 nsew signal output
rlabel metal2 s 70306 199200 70362 200000 6 uP_instr[15]
port 611 nsew signal output
rlabel metal2 s 48226 199200 48282 200000 6 uP_instr[1]
port 612 nsew signal output
rlabel metal2 s 50066 199200 50122 200000 6 uP_instr[2]
port 613 nsew signal output
rlabel metal2 s 51906 199200 51962 200000 6 uP_instr[3]
port 614 nsew signal output
rlabel metal2 s 53746 199200 53802 200000 6 uP_instr[4]
port 615 nsew signal output
rlabel metal2 s 55586 199200 55642 200000 6 uP_instr[5]
port 616 nsew signal output
rlabel metal2 s 57426 199200 57482 200000 6 uP_instr[6]
port 617 nsew signal output
rlabel metal2 s 59266 199200 59322 200000 6 uP_instr[7]
port 618 nsew signal output
rlabel metal2 s 60738 199200 60794 200000 6 uP_instr[8]
port 619 nsew signal output
rlabel metal2 s 62210 199200 62266 200000 6 uP_instr[9]
port 620 nsew signal output
rlabel metal2 s 46754 199200 46810 200000 6 uP_instr_mem_addr[0]
port 621 nsew signal input
rlabel metal2 s 64050 199200 64106 200000 6 uP_instr_mem_addr[10]
port 622 nsew signal input
rlabel metal2 s 65522 199200 65578 200000 6 uP_instr_mem_addr[11]
port 623 nsew signal input
rlabel metal2 s 66994 199200 67050 200000 6 uP_instr_mem_addr[12]
port 624 nsew signal input
rlabel metal2 s 48594 199200 48650 200000 6 uP_instr_mem_addr[1]
port 625 nsew signal input
rlabel metal2 s 50434 199200 50490 200000 6 uP_instr_mem_addr[2]
port 626 nsew signal input
rlabel metal2 s 52274 199200 52330 200000 6 uP_instr_mem_addr[3]
port 627 nsew signal input
rlabel metal2 s 54114 199200 54170 200000 6 uP_instr_mem_addr[4]
port 628 nsew signal input
rlabel metal2 s 55954 199200 56010 200000 6 uP_instr_mem_addr[5]
port 629 nsew signal input
rlabel metal2 s 57794 199200 57850 200000 6 uP_instr_mem_addr[6]
port 630 nsew signal input
rlabel metal2 s 59634 199200 59690 200000 6 uP_instr_mem_addr[7]
port 631 nsew signal input
rlabel metal2 s 61106 199200 61162 200000 6 uP_instr_mem_addr[8]
port 632 nsew signal input
rlabel metal2 s 62578 199200 62634 200000 6 uP_instr_mem_addr[9]
port 633 nsew signal input
rlabel metal2 s 47122 199200 47178 200000 6 uP_read_data[0]
port 634 nsew signal output
rlabel metal2 s 64418 199200 64474 200000 6 uP_read_data[10]
port 635 nsew signal output
rlabel metal2 s 65890 199200 65946 200000 6 uP_read_data[11]
port 636 nsew signal output
rlabel metal2 s 67362 199200 67418 200000 6 uP_read_data[12]
port 637 nsew signal output
rlabel metal2 s 68466 199200 68522 200000 6 uP_read_data[13]
port 638 nsew signal output
rlabel metal2 s 69570 199200 69626 200000 6 uP_read_data[14]
port 639 nsew signal output
rlabel metal2 s 70674 199200 70730 200000 6 uP_read_data[15]
port 640 nsew signal output
rlabel metal2 s 48962 199200 49018 200000 6 uP_read_data[1]
port 641 nsew signal output
rlabel metal2 s 50802 199200 50858 200000 6 uP_read_data[2]
port 642 nsew signal output
rlabel metal2 s 52642 199200 52698 200000 6 uP_read_data[3]
port 643 nsew signal output
rlabel metal2 s 54482 199200 54538 200000 6 uP_read_data[4]
port 644 nsew signal output
rlabel metal2 s 56322 199200 56378 200000 6 uP_read_data[5]
port 645 nsew signal output
rlabel metal2 s 58162 199200 58218 200000 6 uP_read_data[6]
port 646 nsew signal output
rlabel metal2 s 60002 199200 60058 200000 6 uP_read_data[7]
port 647 nsew signal output
rlabel metal2 s 61474 199200 61530 200000 6 uP_read_data[8]
port 648 nsew signal output
rlabel metal2 s 62946 199200 63002 200000 6 uP_read_data[9]
port 649 nsew signal output
rlabel metal2 s 47490 199200 47546 200000 6 uP_write_data[0]
port 650 nsew signal input
rlabel metal2 s 64786 199200 64842 200000 6 uP_write_data[10]
port 651 nsew signal input
rlabel metal2 s 66258 199200 66314 200000 6 uP_write_data[11]
port 652 nsew signal input
rlabel metal2 s 67730 199200 67786 200000 6 uP_write_data[12]
port 653 nsew signal input
rlabel metal2 s 68834 199200 68890 200000 6 uP_write_data[13]
port 654 nsew signal input
rlabel metal2 s 69938 199200 69994 200000 6 uP_write_data[14]
port 655 nsew signal input
rlabel metal2 s 71042 199200 71098 200000 6 uP_write_data[15]
port 656 nsew signal input
rlabel metal2 s 49330 199200 49386 200000 6 uP_write_data[1]
port 657 nsew signal input
rlabel metal2 s 51170 199200 51226 200000 6 uP_write_data[2]
port 658 nsew signal input
rlabel metal2 s 53010 199200 53066 200000 6 uP_write_data[3]
port 659 nsew signal input
rlabel metal2 s 54850 199200 54906 200000 6 uP_write_data[4]
port 660 nsew signal input
rlabel metal2 s 56690 199200 56746 200000 6 uP_write_data[5]
port 661 nsew signal input
rlabel metal2 s 58530 199200 58586 200000 6 uP_write_data[6]
port 662 nsew signal input
rlabel metal2 s 60370 199200 60426 200000 6 uP_write_data[7]
port 663 nsew signal input
rlabel metal2 s 61842 199200 61898 200000 6 uP_write_data[8]
port 664 nsew signal input
rlabel metal2 s 63314 199200 63370 200000 6 uP_write_data[9]
port 665 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 667 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 667 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 667 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 667 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 667 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 667 nsew ground bidirectional
rlabel metal2 s 1950 0 2006 800 6 wb_clk_i
port 668 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wb_rst_i
port 669 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15589642
string GDS_FILE /home/radhe/mpw8/caravel_user_project/openlane/io_interface/runs/23_01_01_02_26/results/signoff/io_interface.magic.gds
string GDS_START 580240
<< end >>

