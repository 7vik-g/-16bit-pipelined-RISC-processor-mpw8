magic
tech sky130B
magscale 1 2
timestamp 1672521598
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 154114 700612 154120 700664
rect 154172 700652 154178 700664
rect 163498 700652 163504 700664
rect 154172 700624 163504 700652
rect 154172 700612 154178 700624
rect 163498 700612 163504 700624
rect 163556 700612 163562 700664
rect 137830 700544 137836 700596
rect 137888 700584 137894 700596
rect 175918 700584 175924 700596
rect 137888 700556 175924 700584
rect 137888 700544 137894 700556
rect 175918 700544 175924 700556
rect 175976 700544 175982 700596
rect 391198 700544 391204 700596
rect 391256 700584 391262 700596
rect 429838 700584 429844 700596
rect 391256 700556 429844 700584
rect 391256 700544 391262 700556
rect 429838 700544 429844 700556
rect 429896 700544 429902 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 191098 700516 191104 700528
rect 105504 700488 191104 700516
rect 105504 700476 105510 700488
rect 191098 700476 191104 700488
rect 191156 700476 191162 700528
rect 410518 700476 410524 700528
rect 410576 700516 410582 700528
rect 494790 700516 494796 700528
rect 410576 700488 494796 700516
rect 410576 700476 410582 700488
rect 494790 700476 494796 700488
rect 494848 700476 494854 700528
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 180058 700448 180064 700460
rect 89220 700420 180064 700448
rect 89220 700408 89226 700420
rect 180058 700408 180064 700420
rect 180116 700408 180122 700460
rect 202138 700408 202144 700460
rect 202196 700448 202202 700460
rect 235166 700448 235172 700460
rect 202196 700420 235172 700448
rect 202196 700408 202202 700420
rect 235166 700408 235172 700420
rect 235224 700408 235230 700460
rect 393958 700408 393964 700460
rect 394016 700448 394022 700460
rect 478506 700448 478512 700460
rect 394016 700420 478512 700448
rect 394016 700408 394022 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 166258 700380 166264 700392
rect 24360 700352 166264 700380
rect 24360 700340 24366 700352
rect 166258 700340 166264 700352
rect 166316 700340 166322 700392
rect 202230 700340 202236 700392
rect 202288 700380 202294 700392
rect 267642 700380 267648 700392
rect 202288 700352 267648 700380
rect 202288 700340 202294 700352
rect 267642 700340 267648 700352
rect 267700 700340 267706 700392
rect 392578 700340 392584 700392
rect 392636 700380 392642 700392
rect 527174 700380 527180 700392
rect 392636 700352 527180 700380
rect 392636 700340 392642 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 192478 700312 192484 700324
rect 40552 700284 192484 700312
rect 40552 700272 40558 700284
rect 192478 700272 192484 700284
rect 192536 700272 192542 700324
rect 202046 700272 202052 700324
rect 202104 700312 202110 700324
rect 283834 700312 283840 700324
rect 202104 700284 283840 700312
rect 202104 700272 202110 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 389818 700272 389824 700324
rect 389876 700312 389882 700324
rect 397454 700312 397460 700324
rect 389876 700284 397460 700312
rect 389876 700272 389882 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 400858 700272 400864 700324
rect 400916 700312 400922 700324
rect 559650 700312 559656 700324
rect 400916 700284 559656 700312
rect 400916 700272 400922 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 8110 700204 8116 700256
rect 8168 700244 8174 700256
rect 14458 700244 14464 700256
rect 8168 700216 14464 700244
rect 8168 700204 8174 700216
rect 14458 700204 14464 700216
rect 14516 700204 14522 700256
rect 407758 699660 407764 699712
rect 407816 699700 407822 699712
rect 413646 699700 413652 699712
rect 407816 699672 413652 699700
rect 407816 699660 407822 699672
rect 413646 699660 413652 699672
rect 413704 699660 413710 699712
rect 382918 696940 382924 696992
rect 382976 696980 382982 696992
rect 580166 696980 580172 696992
rect 382976 696952 580172 696980
rect 382976 696940 382982 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 174538 683176 174544 683188
rect 3476 683148 174544 683176
rect 3476 683136 3482 683148
rect 174538 683136 174544 683148
rect 174596 683136 174602 683188
rect 385678 683136 385684 683188
rect 385736 683176 385742 683188
rect 580166 683176 580172 683188
rect 385736 683148 580172 683176
rect 385736 683136 385742 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 317414 682660 317420 682712
rect 317472 682700 317478 682712
rect 377766 682700 377772 682712
rect 317472 682672 377772 682700
rect 317472 682660 317478 682672
rect 377766 682660 377772 682672
rect 377824 682660 377830 682712
rect 199930 682592 199936 682644
rect 199988 682632 199994 682644
rect 221734 682632 221740 682644
rect 199988 682604 221740 682632
rect 199988 682592 199994 682604
rect 221734 682592 221740 682604
rect 221792 682592 221798 682644
rect 334158 682592 334164 682644
rect 334216 682632 334222 682644
rect 379698 682632 379704 682644
rect 334216 682604 379704 682632
rect 334216 682592 334222 682604
rect 379698 682592 379704 682604
rect 379756 682592 379762 682644
rect 196618 682524 196624 682576
rect 196676 682564 196682 682576
rect 255222 682564 255228 682576
rect 196676 682536 255228 682564
rect 196676 682524 196682 682536
rect 255222 682524 255228 682536
rect 255280 682524 255286 682576
rect 336550 682524 336556 682576
rect 336608 682564 336614 682576
rect 381170 682564 381176 682576
rect 336608 682536 381176 682564
rect 336608 682524 336614 682536
rect 381170 682524 381176 682536
rect 381228 682524 381234 682576
rect 196526 682456 196532 682508
rect 196584 682496 196590 682508
rect 276750 682496 276756 682508
rect 196584 682468 276756 682496
rect 196584 682456 196590 682468
rect 276750 682456 276756 682468
rect 276808 682456 276814 682508
rect 322198 682456 322204 682508
rect 322256 682496 322262 682508
rect 379606 682496 379612 682508
rect 322256 682468 379612 682496
rect 322256 682456 322262 682468
rect 379606 682456 379612 682468
rect 379664 682456 379670 682508
rect 195054 682388 195060 682440
rect 195112 682428 195118 682440
rect 279142 682428 279148 682440
rect 195112 682400 279148 682428
rect 195112 682388 195118 682400
rect 279142 682388 279148 682400
rect 279200 682388 279206 682440
rect 355686 682388 355692 682440
rect 355744 682428 355750 682440
rect 378318 682428 378324 682440
rect 355744 682400 378324 682428
rect 355744 682388 355750 682400
rect 378318 682388 378324 682400
rect 378376 682388 378382 682440
rect 196710 682320 196716 682372
rect 196768 682360 196774 682372
rect 281534 682360 281540 682372
rect 196768 682332 281540 682360
rect 196768 682320 196774 682332
rect 281534 682320 281540 682332
rect 281592 682320 281598 682372
rect 362862 682320 362868 682372
rect 362920 682360 362926 682372
rect 378502 682360 378508 682372
rect 362920 682332 378508 682360
rect 362920 682320 362926 682332
rect 378502 682320 378508 682332
rect 378560 682320 378566 682372
rect 199654 682252 199660 682304
rect 199712 682292 199718 682304
rect 226518 682292 226524 682304
rect 199712 682264 226524 682292
rect 199712 682252 199718 682264
rect 226518 682252 226524 682264
rect 226576 682252 226582 682304
rect 353294 682252 353300 682304
rect 353352 682292 353358 682304
rect 378226 682292 378232 682304
rect 353352 682264 378232 682292
rect 353352 682252 353358 682264
rect 378226 682252 378232 682264
rect 378284 682252 378290 682304
rect 199838 682184 199844 682236
rect 199896 682224 199902 682236
rect 231302 682224 231308 682236
rect 199896 682196 231308 682224
rect 199896 682184 199902 682196
rect 231302 682184 231308 682196
rect 231360 682184 231366 682236
rect 350902 682184 350908 682236
rect 350960 682224 350966 682236
rect 381078 682224 381084 682236
rect 350960 682196 381084 682224
rect 350960 682184 350966 682196
rect 381078 682184 381084 682196
rect 381136 682184 381142 682236
rect 201954 682116 201960 682168
rect 202012 682156 202018 682168
rect 236086 682156 236092 682168
rect 202012 682128 236092 682156
rect 202012 682116 202018 682128
rect 236086 682116 236092 682128
rect 236144 682116 236150 682168
rect 348510 682116 348516 682168
rect 348568 682156 348574 682168
rect 380986 682156 380992 682168
rect 348568 682128 380992 682156
rect 348568 682116 348574 682128
rect 380986 682116 380992 682128
rect 381044 682116 381050 682168
rect 199378 682048 199384 682100
rect 199436 682088 199442 682100
rect 233694 682088 233700 682100
rect 199436 682060 233700 682088
rect 199436 682048 199442 682060
rect 233694 682048 233700 682060
rect 233752 682048 233758 682100
rect 343726 682048 343732 682100
rect 343784 682088 343790 682100
rect 377582 682088 377588 682100
rect 343784 682060 377588 682088
rect 343784 682048 343790 682060
rect 377582 682048 377588 682060
rect 377640 682048 377646 682100
rect 195882 681980 195888 682032
rect 195940 682020 195946 682032
rect 252830 682020 252836 682032
rect 195940 681992 252836 682020
rect 195940 681980 195946 681992
rect 252830 681980 252836 681992
rect 252888 681980 252894 682032
rect 346118 681980 346124 682032
rect 346176 682020 346182 682032
rect 379514 682020 379520 682032
rect 346176 681992 379520 682020
rect 346176 681980 346182 681992
rect 379514 681980 379520 681992
rect 379572 681980 379578 682032
rect 199562 681912 199568 681964
rect 199620 681952 199626 681964
rect 212166 681952 212172 681964
rect 199620 681924 212172 681952
rect 199620 681912 199626 681924
rect 212166 681912 212172 681924
rect 212224 681912 212230 681964
rect 365254 681912 365260 681964
rect 365312 681952 365318 681964
rect 381262 681952 381268 681964
rect 365312 681924 381268 681952
rect 365312 681912 365318 681924
rect 381262 681912 381268 681924
rect 381320 681912 381326 681964
rect 199746 681844 199752 681896
rect 199804 681884 199810 681896
rect 216950 681884 216956 681896
rect 199804 681856 216956 681884
rect 199804 681844 199810 681856
rect 216950 681844 216956 681856
rect 217008 681844 217014 681896
rect 360470 681844 360476 681896
rect 360528 681884 360534 681896
rect 377674 681884 377680 681896
rect 360528 681856 377680 681884
rect 360528 681844 360534 681856
rect 377674 681844 377680 681856
rect 377732 681844 377738 681896
rect 198642 681776 198648 681828
rect 198700 681816 198706 681828
rect 219342 681816 219348 681828
rect 198700 681788 219348 681816
rect 198700 681776 198706 681788
rect 219342 681776 219348 681788
rect 219400 681776 219406 681828
rect 358078 681776 358084 681828
rect 358136 681816 358142 681828
rect 378410 681816 378416 681828
rect 358136 681788 378416 681816
rect 358136 681776 358142 681788
rect 378410 681776 378416 681788
rect 378468 681776 378474 681828
rect 200022 681708 200028 681760
rect 200080 681748 200086 681760
rect 207382 681748 207388 681760
rect 200080 681720 207388 681748
rect 200080 681708 200086 681720
rect 207382 681708 207388 681720
rect 207440 681708 207446 681760
rect 377214 681708 377220 681760
rect 377272 681748 377278 681760
rect 389266 681748 389272 681760
rect 377272 681720 389272 681748
rect 377272 681708 377278 681720
rect 389266 681708 389272 681720
rect 389324 681708 389330 681760
rect 195514 680892 195520 680944
rect 195572 680932 195578 680944
rect 257614 680932 257620 680944
rect 195572 680904 257620 680932
rect 195572 680892 195578 680904
rect 257614 680892 257620 680904
rect 257672 680892 257678 680944
rect 197078 680824 197084 680876
rect 197136 680864 197142 680876
rect 262398 680864 262404 680876
rect 197136 680836 262404 680864
rect 197136 680824 197142 680836
rect 262398 680824 262404 680836
rect 262456 680824 262462 680876
rect 197170 680756 197176 680808
rect 197228 680796 197234 680808
rect 267182 680796 267188 680808
rect 197228 680768 267188 680796
rect 197228 680756 197234 680768
rect 267182 680756 267188 680768
rect 267240 680756 267246 680808
rect 198458 680688 198464 680740
rect 198516 680728 198522 680740
rect 303062 680728 303068 680740
rect 198516 680700 303068 680728
rect 198516 680688 198522 680700
rect 303062 680688 303068 680700
rect 303120 680688 303126 680740
rect 194410 680620 194416 680672
rect 194468 680660 194474 680672
rect 307846 680660 307852 680672
rect 194468 680632 307852 680660
rect 194468 680620 194474 680632
rect 307846 680620 307852 680632
rect 307904 680620 307910 680672
rect 193030 680552 193036 680604
rect 193088 680592 193094 680604
rect 310238 680592 310244 680604
rect 193088 680564 310244 680592
rect 193088 680552 193094 680564
rect 310238 680552 310244 680564
rect 310296 680552 310302 680604
rect 193122 680484 193128 680536
rect 193180 680524 193186 680536
rect 312630 680524 312636 680536
rect 193180 680496 312636 680524
rect 193180 680484 193186 680496
rect 312630 680484 312636 680496
rect 312688 680484 312694 680536
rect 194502 680416 194508 680468
rect 194560 680456 194566 680468
rect 315022 680456 315028 680468
rect 194560 680428 315028 680456
rect 194560 680416 194566 680428
rect 315022 680416 315028 680428
rect 315080 680416 315086 680468
rect 195422 680348 195428 680400
rect 195480 680388 195486 680400
rect 329374 680388 329380 680400
rect 195480 680360 329380 680388
rect 195480 680348 195486 680360
rect 329374 680348 329380 680360
rect 329432 680348 329438 680400
rect 201678 679804 201684 679856
rect 201736 679844 201742 679856
rect 210970 679844 210976 679856
rect 201736 679816 210976 679844
rect 201736 679804 201742 679816
rect 210970 679804 210976 679816
rect 211028 679804 211034 679856
rect 202506 679736 202512 679788
rect 202564 679776 202570 679788
rect 206002 679776 206008 679788
rect 202564 679748 206008 679776
rect 202564 679736 202570 679748
rect 206002 679736 206008 679748
rect 206060 679736 206066 679788
rect 195946 679680 219434 679708
rect 195146 679600 195152 679652
rect 195204 679640 195210 679652
rect 195946 679640 195974 679680
rect 195204 679612 195974 679640
rect 205606 679612 215294 679640
rect 195204 679600 195210 679612
rect 195698 679532 195704 679584
rect 195756 679572 195762 679584
rect 205606 679572 205634 679612
rect 195756 679544 205634 679572
rect 195756 679532 195762 679544
rect 195606 679464 195612 679516
rect 195664 679504 195670 679516
rect 195664 679476 206324 679504
rect 195664 679464 195670 679476
rect 195790 679396 195796 679448
rect 195848 679436 195854 679448
rect 195848 679408 195974 679436
rect 195848 679396 195854 679408
rect 195946 679368 195974 679408
rect 197262 679396 197268 679448
rect 197320 679436 197326 679448
rect 205634 679436 205640 679448
rect 197320 679408 205640 679436
rect 197320 679396 197326 679408
rect 205634 679396 205640 679408
rect 205692 679396 205698 679448
rect 205818 679396 205824 679448
rect 205876 679396 205882 679448
rect 206002 679396 206008 679448
rect 206060 679396 206066 679448
rect 206296 679436 206324 679476
rect 211108 679464 211114 679516
rect 211166 679504 211172 679516
rect 214190 679504 214196 679516
rect 211166 679476 214196 679504
rect 211166 679464 211172 679476
rect 214190 679464 214196 679476
rect 214248 679464 214254 679516
rect 215266 679504 215294 679612
rect 219406 679572 219434 679680
rect 259638 679572 259644 679584
rect 219406 679544 259644 679572
rect 259638 679532 259644 679544
rect 259696 679532 259702 679584
rect 223758 679504 223764 679516
rect 215266 679476 223764 679504
rect 223758 679464 223764 679476
rect 223816 679464 223822 679516
rect 247678 679504 247684 679516
rect 243372 679476 247684 679504
rect 228542 679436 228548 679448
rect 206296 679408 228548 679436
rect 228542 679396 228548 679408
rect 228600 679396 228606 679448
rect 240502 679436 240508 679448
rect 229066 679408 240508 679436
rect 202506 679368 202512 679380
rect 195946 679340 202512 679368
rect 202506 679328 202512 679340
rect 202564 679328 202570 679380
rect 198550 679260 198556 679312
rect 198608 679300 198614 679312
rect 201770 679300 201776 679312
rect 198608 679272 201776 679300
rect 198608 679260 198614 679272
rect 201770 679260 201776 679272
rect 201828 679260 201834 679312
rect 205836 679300 205864 679396
rect 206020 679368 206048 679396
rect 229066 679368 229094 679408
rect 240502 679396 240508 679408
rect 240560 679396 240566 679448
rect 242894 679396 242900 679448
rect 242952 679396 242958 679448
rect 206020 679340 229094 679368
rect 242912 679300 242940 679396
rect 205836 679272 242940 679300
rect 201586 679192 201592 679244
rect 201644 679232 201650 679244
rect 202322 679232 202328 679244
rect 201644 679204 202328 679232
rect 201644 679192 201650 679204
rect 202322 679192 202328 679204
rect 202380 679192 202386 679244
rect 243372 679232 243400 679476
rect 247678 679464 247684 679476
rect 247736 679464 247742 679516
rect 245562 679396 245568 679448
rect 245620 679396 245626 679448
rect 250070 679436 250076 679448
rect 248386 679408 250076 679436
rect 205652 679204 243400 679232
rect 201310 679124 201316 679176
rect 201368 679164 201374 679176
rect 205652 679164 205680 679204
rect 245580 679164 245608 679396
rect 201368 679136 205680 679164
rect 205836 679136 245608 679164
rect 201368 679124 201374 679136
rect 201402 678988 201408 679040
rect 201460 679028 201466 679040
rect 201678 679028 201684 679040
rect 201460 679000 201684 679028
rect 201460 678988 201466 679000
rect 201678 678988 201684 679000
rect 201736 678988 201742 679040
rect 201770 678852 201776 678904
rect 201828 678892 201834 678904
rect 205836 678892 205864 679136
rect 248386 679096 248414 679408
rect 250070 679396 250076 679408
rect 250128 679396 250134 679448
rect 324866 679396 324872 679448
rect 324924 679396 324930 679448
rect 215266 679068 248414 679096
rect 215266 679028 215294 679068
rect 201828 678864 205864 678892
rect 211126 679000 215294 679028
rect 324884 679028 324912 679396
rect 379790 679028 379796 679040
rect 324884 679000 379796 679028
rect 201828 678852 201834 678864
rect 202322 678784 202328 678836
rect 202380 678824 202386 678836
rect 211126 678824 211154 679000
rect 379790 678988 379796 679000
rect 379848 678988 379854 679040
rect 202380 678796 211154 678824
rect 202380 678784 202386 678796
rect 201954 678308 201960 678360
rect 202012 678348 202018 678360
rect 202414 678348 202420 678360
rect 202012 678320 202420 678348
rect 202012 678308 202018 678320
rect 202414 678308 202420 678320
rect 202472 678308 202478 678360
rect 150986 674840 150992 674892
rect 151044 674880 151050 674892
rect 157334 674880 157340 674892
rect 151044 674852 157340 674880
rect 151044 674840 151050 674852
rect 157334 674840 157340 674852
rect 157392 674840 157398 674892
rect 551002 674840 551008 674892
rect 551060 674880 551066 674892
rect 557534 674880 557540 674892
rect 551060 674852 557540 674880
rect 551060 674840 551066 674852
rect 557534 674840 557540 674852
rect 557592 674840 557598 674892
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 10318 670732 10324 670744
rect 3568 670704 10324 670732
rect 3568 670692 3574 670704
rect 10318 670692 10324 670704
rect 10376 670692 10382 670744
rect 565078 670692 565084 670744
rect 565136 670732 565142 670744
rect 580166 670732 580172 670744
rect 565136 670704 580172 670732
rect 565136 670692 565142 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 658112 3424 658164
rect 3476 658152 3482 658164
rect 7558 658152 7564 658164
rect 3476 658124 7564 658152
rect 3476 658112 3482 658124
rect 7558 658112 7564 658124
rect 7616 658112 7622 658164
rect 569218 643084 569224 643136
rect 569276 643124 569282 643136
rect 580166 643124 580172 643136
rect 569276 643096 580172 643124
rect 569276 643084 569282 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 573358 630640 573364 630692
rect 573416 630680 573422 630692
rect 580166 630680 580172 630692
rect 573416 630652 580172 630680
rect 573416 630640 573422 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 14550 618304 14556 618316
rect 3200 618276 14556 618304
rect 3200 618264 3206 618276
rect 14550 618264 14556 618276
rect 14608 618264 14614 618316
rect 563698 616836 563704 616888
rect 563756 616876 563762 616888
rect 580166 616876 580172 616888
rect 563756 616848 580172 616876
rect 563756 616836 563762 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 11698 605860 11704 605872
rect 3292 605832 11704 605860
rect 3292 605820 3298 605832
rect 11698 605820 11704 605832
rect 11756 605820 11762 605872
rect 403618 597524 403624 597576
rect 403676 597564 403682 597576
rect 416774 597564 416780 597576
rect 403676 597536 416780 597564
rect 403676 597524 403682 597536
rect 416774 597524 416780 597536
rect 416832 597524 416838 597576
rect 417786 591336 417792 591388
rect 417844 591376 417850 591388
rect 419442 591376 419448 591388
rect 417844 591348 419448 591376
rect 417844 591336 417850 591348
rect 419442 591336 419448 591348
rect 419500 591336 419506 591388
rect 558178 590656 558184 590708
rect 558236 590696 558242 590708
rect 579798 590696 579804 590708
rect 558236 590668 579804 590696
rect 558236 590656 558242 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 16298 589228 16304 589280
rect 16356 589268 16362 589280
rect 19242 589268 19248 589280
rect 16356 589240 19248 589268
rect 16356 589228 16362 589240
rect 19242 589228 19248 589240
rect 19300 589228 19306 589280
rect 51074 587800 51080 587852
rect 51132 587840 51138 587852
rect 69750 587840 69756 587852
rect 51132 587812 69756 587840
rect 51132 587800 51138 587812
rect 69750 587800 69756 587812
rect 69808 587800 69814 587852
rect 473262 587800 473268 587852
rect 473320 587840 473326 587852
rect 476942 587840 476948 587852
rect 473320 587812 476948 587840
rect 473320 587800 473326 587812
rect 476942 587800 476948 587812
rect 477000 587800 477006 587852
rect 522390 587800 522396 587852
rect 522448 587840 522454 587852
rect 525886 587840 525892 587852
rect 522448 587812 525892 587840
rect 522448 587800 522454 587812
rect 525886 587800 525892 587812
rect 525944 587800 525950 587852
rect 44174 587732 44180 587784
rect 44232 587772 44238 587784
rect 62758 587772 62764 587784
rect 44232 587744 62764 587772
rect 44232 587732 44238 587744
rect 62758 587732 62764 587744
rect 62816 587732 62822 587784
rect 50062 587664 50068 587716
rect 50120 587704 50126 587716
rect 68646 587704 68652 587716
rect 50120 587676 68652 587704
rect 50120 587664 50126 587676
rect 68646 587664 68652 587676
rect 68704 587664 68710 587716
rect 18598 587596 18604 587648
rect 18656 587636 18662 587648
rect 53834 587636 53840 587648
rect 18656 587608 53840 587636
rect 18656 587596 18662 587608
rect 53834 587596 53840 587608
rect 53892 587596 53898 587648
rect 55674 587596 55680 587648
rect 55732 587636 55738 587648
rect 74350 587636 74356 587648
rect 55732 587608 74356 587636
rect 55732 587596 55738 587608
rect 74350 587596 74356 587608
rect 74408 587596 74414 587648
rect 42794 587528 42800 587580
rect 42852 587568 42858 587580
rect 61286 587568 61292 587580
rect 42852 587540 61292 587568
rect 42852 587528 42858 587540
rect 61286 587528 61292 587540
rect 61344 587528 61350 587580
rect 414658 587528 414664 587580
rect 414716 587568 414722 587580
rect 456058 587568 456064 587580
rect 414716 587540 456064 587568
rect 414716 587528 414722 587540
rect 456058 587528 456064 587540
rect 456116 587528 456122 587580
rect 17126 587460 17132 587512
rect 17184 587500 17190 587512
rect 60550 587500 60556 587512
rect 17184 587472 60556 587500
rect 17184 587460 17190 587472
rect 60550 587460 60556 587472
rect 60608 587500 60614 587512
rect 79134 587500 79140 587512
rect 60608 587472 79140 587500
rect 60608 587460 60614 587472
rect 79134 587460 79140 587472
rect 79192 587460 79198 587512
rect 419994 587460 420000 587512
rect 420052 587500 420058 587512
rect 459738 587500 459744 587512
rect 420052 587472 459744 587500
rect 420052 587460 420058 587472
rect 459738 587460 459744 587472
rect 459796 587460 459802 587512
rect 48130 587392 48136 587444
rect 48188 587432 48194 587444
rect 66254 587432 66260 587444
rect 48188 587404 66260 587432
rect 48188 587392 48194 587404
rect 66254 587392 66260 587404
rect 66312 587392 66318 587444
rect 125962 587392 125968 587444
rect 126020 587432 126026 587444
rect 156690 587432 156696 587444
rect 126020 587404 156696 587432
rect 126020 587392 126026 587404
rect 156690 587392 156696 587404
rect 156748 587392 156754 587444
rect 461578 587432 461584 587444
rect 451246 587404 461584 587432
rect 18414 587324 18420 587376
rect 18472 587364 18478 587376
rect 39574 587364 39580 587376
rect 18472 587336 39580 587364
rect 18472 587324 18478 587336
rect 39574 587324 39580 587336
rect 39632 587324 39638 587376
rect 46842 587324 46848 587376
rect 46900 587364 46906 587376
rect 64966 587364 64972 587376
rect 46900 587336 64972 587364
rect 46900 587324 46906 587336
rect 64966 587324 64972 587336
rect 65024 587324 65030 587376
rect 111242 587324 111248 587376
rect 111300 587364 111306 587376
rect 162118 587364 162124 587376
rect 111300 587336 162124 587364
rect 111300 587324 111306 587336
rect 162118 587324 162124 587336
rect 162176 587324 162182 587376
rect 451246 587364 451274 587404
rect 461578 587392 461584 587404
rect 461636 587392 461642 587444
rect 445312 587336 451274 587364
rect 19794 587256 19800 587308
rect 19852 587296 19858 587308
rect 42794 587296 42800 587308
rect 19852 587268 42800 587296
rect 19852 587256 19858 587268
rect 42794 587256 42800 587268
rect 42852 587256 42858 587308
rect 63862 587296 63868 587308
rect 45526 587268 63868 587296
rect 16114 587188 16120 587240
rect 16172 587228 16178 587240
rect 45278 587228 45284 587240
rect 16172 587200 45284 587228
rect 16172 587188 16178 587200
rect 45278 587188 45284 587200
rect 45336 587228 45342 587240
rect 45526 587228 45554 587268
rect 63862 587256 63868 587268
rect 63920 587256 63926 587308
rect 103606 587256 103612 587308
rect 103664 587296 103670 587308
rect 156598 587296 156604 587308
rect 103664 587268 156604 587296
rect 103664 587256 103670 587268
rect 156598 587256 156604 587268
rect 156656 587256 156662 587308
rect 419902 587256 419908 587308
rect 419960 587296 419966 587308
rect 438118 587296 438124 587308
rect 419960 587268 438124 587296
rect 419960 587256 419966 587268
rect 438118 587256 438124 587268
rect 438176 587256 438182 587308
rect 45336 587200 45554 587228
rect 45336 587188 45342 587200
rect 53834 587188 53840 587240
rect 53892 587228 53898 587240
rect 73246 587228 73252 587240
rect 53892 587200 73252 587228
rect 53892 587188 53898 587200
rect 73246 587188 73252 587200
rect 73304 587188 73310 587240
rect 100938 587188 100944 587240
rect 100996 587228 101002 587240
rect 156782 587228 156788 587240
rect 100996 587200 156788 587228
rect 100996 587188 101002 587200
rect 156782 587188 156788 587200
rect 156840 587188 156846 587240
rect 419810 587188 419816 587240
rect 419868 587228 419874 587240
rect 439590 587228 439596 587240
rect 419868 587200 439596 587228
rect 419868 587188 419874 587200
rect 439590 587188 439596 587200
rect 439648 587188 439654 587240
rect 19978 587120 19984 587172
rect 20036 587160 20042 587172
rect 48590 587160 48596 587172
rect 20036 587132 48596 587160
rect 20036 587120 20042 587132
rect 48590 587120 48596 587132
rect 48648 587160 48654 587172
rect 67634 587160 67640 587172
rect 48648 587132 67640 587160
rect 48648 587120 48654 587132
rect 67634 587120 67640 587132
rect 67692 587120 67698 587172
rect 98546 587120 98552 587172
rect 98604 587160 98610 587172
rect 158070 587160 158076 587172
rect 98604 587132 158076 587160
rect 98604 587120 98610 587132
rect 158070 587120 158076 587132
rect 158128 587120 158134 587172
rect 417694 587120 417700 587172
rect 417752 587160 417758 587172
rect 441614 587160 441620 587172
rect 417752 587132 441620 587160
rect 417752 587120 417758 587132
rect 441614 587120 441620 587132
rect 441672 587120 441678 587172
rect 16390 587052 16396 587104
rect 16448 587092 16454 587104
rect 46842 587092 46848 587104
rect 16448 587064 46848 587092
rect 16448 587052 16454 587064
rect 46842 587052 46848 587064
rect 46900 587052 46906 587104
rect 96062 587052 96068 587104
rect 96120 587092 96126 587104
rect 159450 587092 159456 587104
rect 96120 587064 159456 587092
rect 96120 587052 96126 587064
rect 159450 587052 159456 587064
rect 159508 587052 159514 587104
rect 413922 587052 413928 587104
rect 413980 587092 413986 587104
rect 443086 587092 443092 587104
rect 413980 587064 443092 587092
rect 413980 587052 413986 587064
rect 443086 587052 443092 587064
rect 443144 587092 443150 587104
rect 445312 587092 445340 587336
rect 452654 587324 452660 587376
rect 452712 587364 452718 587376
rect 454586 587364 454592 587376
rect 452712 587336 454592 587364
rect 452712 587324 452718 587336
rect 454586 587324 454592 587336
rect 454644 587364 454650 587376
rect 473354 587364 473360 587376
rect 454644 587336 473360 587364
rect 454644 587324 454650 587336
rect 473354 587324 473360 587336
rect 473412 587324 473418 587376
rect 445662 587256 445668 587308
rect 445720 587296 445726 587308
rect 463878 587296 463884 587308
rect 445720 587268 463884 587296
rect 445720 587256 445726 587268
rect 463878 587256 463884 587268
rect 463936 587256 463942 587308
rect 462774 587228 462780 587240
rect 443144 587064 445340 587092
rect 445404 587200 462780 587228
rect 443144 587052 443150 587064
rect 15102 586984 15108 587036
rect 15160 587024 15166 587036
rect 44174 587024 44180 587036
rect 15160 586996 44180 587024
rect 15160 586984 15166 586996
rect 44174 586984 44180 586996
rect 44232 586984 44238 587036
rect 93578 586984 93584 587036
rect 93636 587024 93642 587036
rect 158162 587024 158168 587036
rect 93636 586996 158168 587024
rect 93636 586984 93642 586996
rect 158162 586984 158168 586996
rect 158220 586984 158226 587036
rect 413738 586984 413744 587036
rect 413796 587024 413802 587036
rect 444190 587024 444196 587036
rect 413796 586996 444196 587024
rect 413796 586984 413802 586996
rect 444190 586984 444196 586996
rect 444248 587024 444254 587036
rect 445404 587024 445432 587200
rect 462774 587188 462780 587200
rect 462832 587188 462838 587240
rect 449894 587120 449900 587172
rect 449952 587160 449958 587172
rect 450814 587160 450820 587172
rect 449952 587132 450820 587160
rect 449952 587120 449958 587132
rect 450814 587120 450820 587132
rect 450872 587120 450878 587172
rect 459738 587120 459744 587172
rect 459796 587160 459802 587172
rect 460658 587160 460664 587172
rect 459796 587132 460664 587160
rect 459796 587120 459802 587132
rect 460658 587120 460664 587132
rect 460716 587160 460722 587172
rect 479150 587160 479156 587172
rect 460716 587132 479156 587160
rect 460716 587120 460722 587132
rect 479150 587120 479156 587132
rect 479208 587120 479214 587172
rect 448514 587052 448520 587104
rect 448572 587092 448578 587104
rect 467558 587092 467564 587104
rect 448572 587064 467564 587092
rect 448572 587052 448578 587064
rect 467558 587052 467564 587064
rect 467616 587052 467622 587104
rect 450630 587024 450636 587036
rect 444248 586996 445432 587024
rect 449820 586996 450636 587024
rect 444248 586984 444254 586996
rect 19702 586916 19708 586968
rect 19760 586956 19766 586968
rect 51074 586956 51080 586968
rect 19760 586928 51080 586956
rect 19760 586916 19766 586928
rect 51074 586916 51080 586928
rect 51132 586916 51138 586968
rect 88242 586916 88248 586968
rect 88300 586956 88306 586968
rect 159358 586956 159364 586968
rect 88300 586928 159364 586956
rect 88300 586916 88306 586928
rect 159358 586916 159364 586928
rect 159416 586916 159422 586968
rect 418798 586916 418804 586968
rect 418856 586956 418862 586968
rect 449820 586956 449848 586996
rect 450630 586984 450636 586996
rect 450688 586984 450694 587036
rect 466270 587024 466276 587036
rect 450740 586996 466276 587024
rect 418856 586928 449848 586956
rect 418856 586916 418862 586928
rect 15010 586848 15016 586900
rect 15068 586888 15074 586900
rect 48130 586888 48136 586900
rect 15068 586860 48136 586888
rect 15068 586848 15074 586860
rect 48130 586848 48136 586860
rect 48188 586848 48194 586900
rect 83642 586848 83648 586900
rect 83700 586888 83706 586900
rect 158254 586888 158260 586900
rect 83700 586860 158260 586888
rect 83700 586848 83706 586860
rect 158254 586848 158260 586860
rect 158312 586848 158318 586900
rect 413830 586848 413836 586900
rect 413888 586888 413894 586900
rect 445662 586888 445668 586900
rect 413888 586860 445668 586888
rect 413888 586848 413894 586860
rect 445662 586848 445668 586860
rect 445720 586848 445726 586900
rect 447318 586848 447324 586900
rect 447376 586888 447382 586900
rect 450740 586888 450768 586996
rect 466270 586984 466276 586996
rect 466328 586984 466334 587036
rect 450814 586916 450820 586968
rect 450872 586956 450878 586968
rect 468662 586956 468668 586968
rect 450872 586928 468668 586956
rect 450872 586916 450878 586928
rect 468662 586916 468668 586928
rect 468720 586916 468726 586968
rect 465166 586888 465172 586900
rect 447376 586860 450768 586888
rect 451246 586860 465172 586888
rect 447376 586848 447382 586860
rect 16482 586780 16488 586832
rect 16540 586820 16546 586832
rect 50062 586820 50068 586832
rect 16540 586792 50068 586820
rect 16540 586780 16546 586792
rect 50062 586780 50068 586792
rect 50120 586780 50126 586832
rect 51074 586780 51080 586832
rect 51132 586820 51138 586832
rect 52362 586820 52368 586832
rect 51132 586792 52368 586820
rect 51132 586780 51138 586792
rect 52362 586780 52368 586792
rect 52420 586820 52426 586832
rect 71130 586820 71136 586832
rect 52420 586792 71136 586820
rect 52420 586780 52426 586792
rect 71130 586780 71136 586792
rect 71188 586780 71194 586832
rect 91002 586780 91008 586832
rect 91060 586820 91066 586832
rect 166350 586820 166356 586832
rect 91060 586792 166356 586820
rect 91060 586780 91066 586792
rect 166350 586780 166356 586792
rect 166408 586780 166414 586832
rect 445754 586780 445760 586832
rect 445812 586820 445818 586832
rect 446490 586820 446496 586832
rect 445812 586792 446496 586820
rect 445812 586780 445818 586792
rect 446490 586780 446496 586792
rect 446548 586820 446554 586832
rect 451246 586820 451274 586860
rect 465166 586848 465172 586860
rect 465224 586848 465230 586900
rect 446548 586792 451274 586820
rect 446548 586780 446554 586792
rect 451366 586780 451372 586832
rect 451424 586820 451430 586832
rect 469766 586820 469772 586832
rect 451424 586792 469772 586820
rect 451424 586780 451430 586792
rect 469766 586780 469772 586792
rect 469824 586780 469830 586832
rect 52638 586712 52644 586764
rect 52696 586752 52702 586764
rect 72142 586752 72148 586764
rect 52696 586724 72148 586752
rect 52696 586712 52702 586724
rect 72142 586712 72148 586724
rect 72200 586712 72206 586764
rect 73706 586712 73712 586764
rect 73764 586752 73770 586764
rect 157978 586752 157984 586764
rect 73764 586724 157984 586752
rect 73764 586712 73770 586724
rect 157978 586712 157984 586724
rect 158036 586712 158042 586764
rect 451274 586712 451280 586764
rect 451332 586752 451338 586764
rect 452378 586752 452384 586764
rect 451332 586724 452384 586752
rect 451332 586712 451338 586724
rect 452378 586712 452384 586724
rect 452436 586752 452442 586764
rect 471238 586752 471244 586764
rect 452436 586724 471244 586752
rect 452436 586712 452442 586724
rect 471238 586712 471244 586724
rect 471296 586712 471302 586764
rect 15838 586644 15844 586696
rect 15896 586684 15902 586696
rect 55674 586684 55680 586696
rect 15896 586656 55680 586684
rect 15896 586644 15902 586656
rect 55674 586644 55680 586656
rect 55732 586644 55738 586696
rect 78490 586644 78496 586696
rect 78548 586684 78554 586696
rect 163590 586684 163596 586696
rect 78548 586656 163596 586684
rect 78548 586644 78554 586656
rect 163590 586644 163596 586656
rect 163648 586644 163654 586696
rect 419718 586644 419724 586696
rect 419776 586684 419782 586696
rect 452654 586684 452660 586696
rect 419776 586656 452660 586684
rect 419776 586644 419782 586656
rect 452654 586644 452660 586656
rect 452712 586644 452718 586696
rect 452746 586644 452752 586696
rect 452804 586684 452810 586696
rect 453482 586684 453488 586696
rect 452804 586656 453488 586684
rect 452804 586644 452810 586656
rect 453482 586644 453488 586656
rect 453540 586684 453546 586696
rect 453540 586656 453712 586684
rect 453540 586644 453546 586656
rect 16206 586576 16212 586628
rect 16264 586616 16270 586628
rect 57054 586616 57060 586628
rect 16264 586588 57060 586616
rect 16264 586576 16270 586588
rect 57054 586576 57060 586588
rect 57112 586576 57118 586628
rect 76098 586576 76104 586628
rect 76156 586616 76162 586628
rect 162210 586616 162216 586628
rect 76156 586588 162216 586616
rect 76156 586576 76162 586588
rect 162210 586576 162216 586588
rect 162268 586576 162274 586628
rect 416038 586576 416044 586628
rect 416096 586616 416102 586628
rect 453574 586616 453580 586628
rect 416096 586588 453580 586616
rect 416096 586576 416102 586588
rect 453574 586576 453580 586588
rect 453632 586576 453638 586628
rect 453684 586616 453712 586656
rect 456150 586644 456156 586696
rect 456208 586684 456214 586696
rect 473630 586684 473636 586696
rect 456208 586656 473636 586684
rect 456208 586644 456214 586656
rect 473630 586644 473636 586656
rect 473688 586644 473694 586696
rect 472158 586616 472164 586628
rect 453684 586588 472164 586616
rect 472158 586576 472164 586588
rect 472216 586576 472222 586628
rect 474090 586576 474096 586628
rect 474148 586616 474154 586628
rect 523310 586616 523316 586628
rect 474148 586588 523316 586616
rect 474148 586576 474154 586588
rect 523310 586576 523316 586588
rect 523368 586576 523374 586628
rect 19886 586508 19892 586560
rect 19944 586548 19950 586560
rect 36630 586548 36636 586560
rect 19944 586520 36636 586548
rect 19944 586508 19950 586520
rect 36630 586508 36636 586520
rect 36688 586508 36694 586560
rect 59814 586508 59820 586560
rect 59872 586548 59878 586560
rect 77386 586548 77392 586560
rect 59872 586520 77392 586548
rect 59872 586508 59878 586520
rect 77386 586508 77392 586520
rect 77444 586508 77450 586560
rect 81066 586508 81072 586560
rect 81124 586548 81130 586560
rect 167638 586548 167644 586560
rect 81124 586520 167644 586548
rect 81124 586508 81130 586520
rect 167638 586508 167644 586520
rect 167696 586508 167702 586560
rect 380158 586508 380164 586560
rect 380216 586548 380222 586560
rect 458174 586548 458180 586560
rect 380216 586520 458180 586548
rect 380216 586508 380222 586520
rect 458174 586508 458180 586520
rect 458232 586508 458238 586560
rect 458266 586508 458272 586560
rect 458324 586548 458330 586560
rect 478046 586548 478052 586560
rect 458324 586520 478052 586548
rect 458324 586508 458330 586520
rect 478046 586508 478052 586520
rect 478104 586508 478110 586560
rect 19242 586440 19248 586492
rect 19300 586480 19306 586492
rect 150710 586480 150716 586492
rect 19300 586452 150716 586480
rect 19300 586440 19306 586452
rect 150710 586440 150716 586452
rect 150768 586480 150774 586492
rect 157334 586480 157340 586492
rect 150768 586452 157340 586480
rect 150768 586440 150774 586452
rect 157334 586440 157340 586452
rect 157392 586440 157398 586492
rect 417786 586440 417792 586492
rect 417844 586480 417850 586492
rect 550818 586480 550824 586492
rect 417844 586452 550824 586480
rect 417844 586440 417850 586452
rect 550818 586440 550824 586452
rect 550876 586480 550882 586492
rect 557534 586480 557540 586492
rect 550876 586452 557540 586480
rect 550876 586440 550882 586452
rect 557534 586440 557540 586452
rect 557592 586440 557598 586492
rect 417694 586372 417700 586424
rect 417752 586412 417758 586424
rect 449894 586412 449900 586424
rect 417752 586384 449900 586412
rect 417752 586372 417758 586384
rect 449894 586372 449900 586384
rect 449952 586372 449958 586424
rect 419350 586304 419356 586356
rect 419408 586344 419414 586356
rect 452746 586344 452752 586356
rect 419408 586316 452752 586344
rect 419408 586304 419414 586316
rect 452746 586304 452752 586316
rect 452804 586304 452810 586356
rect 417326 586236 417332 586288
rect 417384 586276 417390 586288
rect 451274 586276 451280 586288
rect 417384 586248 451280 586276
rect 417384 586236 417390 586248
rect 451274 586236 451280 586248
rect 451332 586236 451338 586288
rect 418614 586168 418620 586220
rect 418672 586208 418678 586220
rect 456150 586208 456156 586220
rect 418672 586180 456156 586208
rect 418672 586168 418678 586180
rect 456150 586168 456156 586180
rect 456208 586168 456214 586220
rect 415854 586100 415860 586152
rect 415912 586140 415918 586152
rect 456794 586140 456800 586152
rect 415912 586112 456800 586140
rect 415912 586100 415918 586112
rect 456794 586100 456800 586112
rect 456852 586100 456858 586152
rect 378962 586032 378968 586084
rect 379020 586032 379026 586084
rect 379054 586032 379060 586084
rect 379112 586072 379118 586084
rect 462314 586072 462320 586084
rect 379112 586044 462320 586072
rect 379112 586032 379118 586044
rect 462314 586032 462320 586044
rect 462372 586032 462378 586084
rect 378980 586004 379008 586032
rect 470594 586004 470600 586016
rect 378980 585976 470600 586004
rect 470594 585964 470600 585976
rect 470652 585964 470658 586016
rect 378962 585896 378968 585948
rect 379020 585936 379026 585948
rect 513374 585936 513380 585948
rect 379020 585908 513380 585936
rect 379020 585896 379026 585908
rect 513374 585896 513380 585908
rect 513432 585896 513438 585948
rect 385034 585828 385040 585880
rect 385092 585868 385098 585880
rect 522390 585868 522396 585880
rect 385092 585840 522396 585868
rect 385092 585828 385098 585840
rect 522390 585828 522396 585840
rect 522448 585828 522454 585880
rect 379054 585760 379060 585812
rect 379112 585800 379118 585812
rect 520274 585800 520280 585812
rect 379112 585772 520280 585800
rect 379112 585760 379118 585772
rect 520274 585760 520280 585772
rect 520332 585760 520338 585812
rect 108390 585080 108396 585132
rect 108448 585120 108454 585132
rect 200850 585120 200856 585132
rect 108448 585092 200856 585120
rect 108448 585080 108454 585092
rect 200850 585080 200856 585092
rect 200908 585080 200914 585132
rect 418890 585080 418896 585132
rect 418948 585120 418954 585132
rect 485774 585120 485780 585132
rect 418948 585092 485780 585120
rect 418948 585080 418954 585092
rect 485774 585080 485780 585092
rect 485832 585080 485838 585132
rect 105538 585012 105544 585064
rect 105596 585052 105602 585064
rect 200942 585052 200948 585064
rect 105596 585024 200948 585052
rect 105596 585012 105602 585024
rect 200942 585012 200948 585024
rect 201000 585012 201006 585064
rect 416590 585012 416596 585064
rect 416648 585052 416654 585064
rect 487154 585052 487160 585064
rect 416648 585024 487160 585052
rect 416648 585012 416654 585024
rect 487154 585012 487160 585024
rect 487212 585012 487218 585064
rect 68554 584944 68560 584996
rect 68612 584984 68618 584996
rect 197814 584984 197820 584996
rect 68612 584956 197820 584984
rect 68612 584944 68618 584956
rect 197814 584944 197820 584956
rect 197872 584944 197878 584996
rect 416498 584944 416504 584996
rect 416556 584984 416562 584996
rect 489914 584984 489920 584996
rect 416556 584956 489920 584984
rect 416556 584944 416562 584956
rect 489914 584944 489920 584956
rect 489972 584944 489978 584996
rect 65978 584876 65984 584928
rect 66036 584916 66042 584928
rect 197906 584916 197912 584928
rect 66036 584888 197912 584916
rect 66036 584876 66042 584888
rect 197906 584876 197912 584888
rect 197964 584876 197970 584928
rect 416222 584876 416228 584928
rect 416280 584916 416286 584928
rect 492674 584916 492680 584928
rect 416280 584888 492680 584916
rect 416280 584876 416286 584888
rect 492674 584876 492680 584888
rect 492732 584876 492738 584928
rect 63954 584808 63960 584860
rect 64012 584848 64018 584860
rect 198182 584848 198188 584860
rect 64012 584820 198188 584848
rect 64012 584808 64018 584820
rect 198182 584808 198188 584820
rect 198240 584808 198246 584860
rect 416682 584808 416688 584860
rect 416740 584848 416746 584860
rect 495434 584848 495440 584860
rect 416740 584820 495440 584848
rect 416740 584808 416746 584820
rect 495434 584808 495440 584820
rect 495492 584808 495498 584860
rect 17034 584740 17040 584792
rect 17092 584780 17098 584792
rect 59814 584780 59820 584792
rect 17092 584752 59820 584780
rect 17092 584740 17098 584752
rect 59814 584740 59820 584752
rect 59872 584740 59878 584792
rect 61838 584740 61844 584792
rect 61896 584780 61902 584792
rect 198274 584780 198280 584792
rect 61896 584752 198280 584780
rect 61896 584740 61902 584752
rect 198274 584740 198280 584752
rect 198332 584740 198338 584792
rect 416314 584740 416320 584792
rect 416372 584780 416378 584792
rect 498194 584780 498200 584792
rect 416372 584752 498200 584780
rect 416372 584740 416378 584752
rect 498194 584740 498200 584752
rect 498252 584740 498258 584792
rect 59262 584672 59268 584724
rect 59320 584712 59326 584724
rect 198366 584712 198372 584724
rect 59320 584684 198372 584712
rect 59320 584672 59326 584684
rect 198366 584672 198372 584684
rect 198424 584672 198430 584724
rect 416406 584672 416412 584724
rect 416464 584712 416470 584724
rect 500954 584712 500960 584724
rect 416464 584684 500960 584712
rect 416464 584672 416470 584684
rect 500954 584672 500960 584684
rect 501012 584672 501018 584724
rect 19058 584604 19064 584656
rect 19116 584644 19122 584656
rect 51074 584644 51080 584656
rect 19116 584616 51080 584644
rect 19116 584604 19122 584616
rect 51074 584604 51080 584616
rect 51132 584604 51138 584656
rect 56226 584604 56232 584656
rect 56284 584644 56290 584656
rect 197998 584644 198004 584656
rect 56284 584616 198004 584644
rect 56284 584604 56290 584616
rect 197998 584604 198004 584616
rect 198056 584604 198062 584656
rect 415946 584604 415952 584656
rect 416004 584644 416010 584656
rect 502334 584644 502340 584656
rect 416004 584616 502340 584644
rect 416004 584604 416010 584616
rect 502334 584604 502340 584616
rect 502392 584604 502398 584656
rect 14918 584536 14924 584588
rect 14976 584576 14982 584588
rect 52638 584576 52644 584588
rect 14976 584548 52644 584576
rect 14976 584536 14982 584548
rect 52638 584536 52644 584548
rect 52696 584536 52702 584588
rect 53650 584536 53656 584588
rect 53708 584576 53714 584588
rect 198090 584576 198096 584588
rect 53708 584548 198096 584576
rect 53708 584536 53714 584548
rect 198090 584536 198096 584548
rect 198148 584536 198154 584588
rect 416130 584536 416136 584588
rect 416188 584576 416194 584588
rect 505094 584576 505100 584588
rect 416188 584548 505100 584576
rect 416188 584536 416194 584548
rect 505094 584536 505100 584548
rect 505152 584536 505158 584588
rect 49786 584468 49792 584520
rect 49844 584508 49850 584520
rect 200666 584508 200672 584520
rect 49844 584480 200672 584508
rect 49844 584468 49850 584480
rect 200666 584468 200672 584480
rect 200724 584468 200730 584520
rect 380894 584468 380900 584520
rect 380952 584508 380958 584520
rect 474090 584508 474096 584520
rect 380952 584480 474096 584508
rect 380952 584468 380958 584480
rect 474090 584468 474096 584480
rect 474148 584468 474154 584520
rect 48682 584400 48688 584452
rect 48740 584440 48746 584452
rect 200574 584440 200580 584452
rect 48740 584412 200580 584440
rect 48740 584400 48746 584412
rect 200574 584400 200580 584412
rect 200632 584400 200638 584452
rect 379146 584400 379152 584452
rect 379204 584440 379210 584452
rect 510614 584440 510620 584452
rect 379204 584412 510620 584440
rect 379204 584400 379210 584412
rect 510614 584400 510620 584412
rect 510672 584400 510678 584452
rect 113818 584332 113824 584384
rect 113876 584372 113882 584384
rect 200758 584372 200764 584384
rect 113876 584344 200764 584372
rect 113876 584332 113882 584344
rect 200758 584332 200764 584344
rect 200816 584332 200822 584384
rect 419258 584332 419264 584384
rect 419316 584372 419322 584384
rect 483014 584372 483020 584384
rect 419316 584344 483020 584372
rect 419316 584332 419322 584344
rect 483014 584332 483020 584344
rect 483072 584332 483078 584384
rect 114554 584264 114560 584316
rect 114612 584304 114618 584316
rect 200850 584304 200856 584316
rect 114612 584276 200856 584304
rect 114612 584264 114618 584276
rect 200850 584264 200856 584276
rect 200908 584264 200914 584316
rect 419074 584264 419080 584316
rect 419132 584304 419138 584316
rect 480254 584304 480260 584316
rect 419132 584276 480260 584304
rect 419132 584264 419138 584276
rect 480254 584264 480260 584276
rect 480312 584264 480318 584316
rect 414842 584196 414848 584248
rect 414900 584236 414906 584248
rect 457254 584236 457260 584248
rect 414900 584208 457260 584236
rect 414900 584196 414906 584208
rect 457254 584196 457260 584208
rect 457312 584196 457318 584248
rect 419442 583516 419448 583568
rect 419500 583556 419506 583568
rect 445754 583556 445760 583568
rect 419500 583528 445760 583556
rect 419500 583516 419506 583528
rect 445754 583516 445760 583528
rect 445812 583516 445818 583568
rect 414750 583448 414756 583500
rect 414808 583488 414814 583500
rect 447318 583488 447324 583500
rect 414808 583460 447324 583488
rect 414808 583448 414814 583460
rect 447318 583448 447324 583460
rect 447376 583448 447382 583500
rect 415026 583380 415032 583432
rect 415084 583420 415090 583432
rect 448514 583420 448520 583432
rect 415084 583392 448520 583420
rect 415084 583380 415090 583392
rect 448514 583380 448520 583392
rect 448572 583380 448578 583432
rect 417234 583312 417240 583364
rect 417292 583352 417298 583364
rect 451366 583352 451372 583364
rect 417292 583324 451372 583352
rect 417292 583312 417298 583324
rect 451366 583312 451372 583324
rect 451424 583312 451430 583364
rect 458266 583312 458272 583364
rect 458324 583312 458330 583364
rect 414934 583244 414940 583296
rect 414992 583284 414998 583296
rect 458284 583284 458312 583312
rect 414992 583256 458312 583284
rect 414992 583244 414998 583256
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 10410 579680 10416 579692
rect 3384 579652 10416 579680
rect 3384 579640 3390 579652
rect 10410 579640 10416 579652
rect 10468 579640 10474 579692
rect 571978 576852 571984 576904
rect 572036 576892 572042 576904
rect 580166 576892 580172 576904
rect 572036 576864 580172 576892
rect 572036 576852 572042 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 562318 563048 562324 563100
rect 562376 563088 562382 563100
rect 579798 563088 579804 563100
rect 562376 563060 579804 563088
rect 562376 563048 562382 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553528 3332 553580
rect 3384 553568 3390 553580
rect 7650 553568 7656 553580
rect 3384 553540 7656 553568
rect 3384 553528 3390 553540
rect 7650 553528 7656 553540
rect 7708 553528 7714 553580
rect 406378 537480 406384 537532
rect 406436 537520 406442 537532
rect 417510 537520 417516 537532
rect 406436 537492 417516 537520
rect 406436 537480 406442 537492
rect 417510 537480 417516 537492
rect 417568 537480 417574 537532
rect 566458 536800 566464 536852
rect 566516 536840 566522 536852
rect 580166 536840 580172 536852
rect 566516 536812 580172 536840
rect 566516 536800 566522 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 383010 536052 383016 536104
rect 383068 536092 383074 536104
rect 417142 536092 417148 536104
rect 383068 536064 417148 536092
rect 383068 536052 383074 536064
rect 417142 536052 417148 536064
rect 417200 536052 417206 536104
rect 415854 535508 415860 535560
rect 415912 535548 415918 535560
rect 416774 535548 416780 535560
rect 415912 535520 416780 535548
rect 415912 535508 415918 535520
rect 416774 535508 416780 535520
rect 416832 535508 416838 535560
rect 417878 535440 417884 535492
rect 417936 535480 417942 535492
rect 418614 535480 418620 535492
rect 417936 535452 418620 535480
rect 417936 535440 417942 535452
rect 418614 535440 418620 535452
rect 418672 535440 418678 535492
rect 414566 533672 414572 533724
rect 414624 533712 414630 533724
rect 417510 533712 417516 533724
rect 414624 533684 417516 533712
rect 414624 533672 414630 533684
rect 417510 533672 417516 533684
rect 417568 533672 417574 533724
rect 17402 531224 17408 531276
rect 17460 531264 17466 531276
rect 18782 531264 18788 531276
rect 17460 531236 18788 531264
rect 17460 531224 17466 531236
rect 18782 531224 18788 531236
rect 18840 531224 18846 531276
rect 411898 530612 411904 530664
rect 411956 530652 411962 530664
rect 416866 530652 416872 530664
rect 411956 530624 416872 530652
rect 411956 530612 411962 530624
rect 416866 530612 416872 530624
rect 416924 530612 416930 530664
rect 410610 530544 410616 530596
rect 410668 530584 410674 530596
rect 416958 530584 416964 530596
rect 410668 530556 416964 530584
rect 410668 530544 410674 530556
rect 416958 530544 416964 530556
rect 417016 530584 417022 530596
rect 417602 530584 417608 530596
rect 417016 530556 417608 530584
rect 417016 530544 417022 530556
rect 417602 530544 417608 530556
rect 417660 530544 417666 530596
rect 16758 528572 16764 528624
rect 16816 528612 16822 528624
rect 19334 528612 19340 528624
rect 16816 528584 19340 528612
rect 16816 528572 16822 528584
rect 19334 528572 19340 528584
rect 19392 528572 19398 528624
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 11790 527184 11796 527196
rect 3016 527156 11796 527184
rect 3016 527144 3022 527156
rect 11790 527144 11796 527156
rect 11848 527144 11854 527196
rect 570598 524424 570604 524476
rect 570656 524464 570662 524476
rect 580166 524464 580172 524476
rect 570656 524436 580172 524464
rect 570656 524424 570662 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 16666 523744 16672 523796
rect 16724 523784 16730 523796
rect 18782 523784 18788 523796
rect 16724 523756 18788 523784
rect 16724 523744 16730 523756
rect 18782 523744 18788 523756
rect 18840 523744 18846 523796
rect 16850 523676 16856 523728
rect 16908 523716 16914 523728
rect 17770 523716 17776 523728
rect 16908 523688 17776 523716
rect 16908 523676 16914 523688
rect 17770 523676 17776 523688
rect 17828 523676 17834 523728
rect 558270 510620 558276 510672
rect 558328 510660 558334 510672
rect 580166 510660 580172 510672
rect 558328 510632 580172 510660
rect 558328 510620 558334 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 17310 510552 17316 510604
rect 17368 510592 17374 510604
rect 19242 510592 19248 510604
rect 17368 510564 19248 510592
rect 17368 510552 17374 510564
rect 19242 510552 19248 510564
rect 19300 510552 19306 510604
rect 387058 509872 387064 509924
rect 387116 509912 387122 509924
rect 416866 509912 416872 509924
rect 387116 509884 416872 509912
rect 387116 509872 387122 509884
rect 416866 509872 416872 509884
rect 416924 509872 416930 509924
rect 389910 507832 389916 507884
rect 389968 507872 389974 507884
rect 417786 507872 417792 507884
rect 389968 507844 417792 507872
rect 389968 507832 389974 507844
rect 417786 507832 417792 507844
rect 417844 507832 417850 507884
rect 365686 501384 367094 501412
rect 202046 501304 202052 501356
rect 202104 501344 202110 501356
rect 202104 501316 209774 501344
rect 202104 501304 202110 501316
rect 209746 501276 209774 501316
rect 209746 501248 211154 501276
rect 211126 501072 211154 501248
rect 365686 501208 365714 501384
rect 367066 501344 367094 501384
rect 367066 501316 371234 501344
rect 353266 501180 354674 501208
rect 211356 501112 211660 501140
rect 211356 501072 211384 501112
rect 211126 501044 211384 501072
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 15746 501004 15752 501016
rect 3384 500976 15752 501004
rect 3384 500964 3390 500976
rect 15746 500964 15752 500976
rect 15804 500964 15810 501016
rect 202230 500964 202236 501016
rect 202288 501004 202294 501016
rect 202288 500976 211154 501004
rect 202288 500964 202294 500976
rect 211126 500954 211154 500976
rect 211632 500954 211660 501112
rect 211126 500926 211476 500954
rect 202138 500760 202144 500812
rect 202196 500800 202202 500812
rect 211448 500800 211476 500926
rect 211540 500926 211660 500954
rect 214116 500976 214420 501004
rect 211540 500868 211568 500926
rect 214116 500868 214144 500976
rect 211540 500840 214144 500868
rect 214392 500868 214420 500976
rect 353266 500936 353294 501180
rect 350506 500908 353294 500936
rect 214392 500840 215616 500868
rect 202196 500772 207704 500800
rect 211448 500772 214328 500800
rect 202196 500760 202202 500772
rect 201954 500692 201960 500744
rect 202012 500732 202018 500744
rect 207566 500732 207572 500744
rect 202012 500704 207572 500732
rect 202012 500692 202018 500704
rect 207566 500692 207572 500704
rect 207624 500692 207630 500744
rect 207676 500732 207704 500772
rect 214300 500744 214328 500772
rect 215588 500744 215616 500840
rect 350506 500800 350534 500908
rect 349356 500772 350534 500800
rect 349356 500744 349384 500772
rect 213362 500732 213368 500744
rect 207676 500704 213368 500732
rect 213362 500692 213368 500704
rect 213420 500692 213426 500744
rect 214282 500692 214288 500744
rect 214340 500692 214346 500744
rect 215570 500692 215576 500744
rect 215628 500692 215634 500744
rect 215662 500692 215668 500744
rect 215720 500732 215726 500744
rect 228358 500732 228364 500744
rect 215720 500704 228364 500732
rect 215720 500692 215726 500704
rect 228358 500692 228364 500704
rect 228416 500692 228422 500744
rect 349338 500692 349344 500744
rect 349396 500692 349402 500744
rect 351822 500732 351828 500744
rect 349448 500704 351828 500732
rect 175918 500624 175924 500676
rect 175976 500664 175982 500676
rect 216950 500664 216956 500676
rect 175976 500636 216956 500664
rect 175976 500624 175982 500636
rect 216950 500624 216956 500636
rect 217008 500624 217014 500676
rect 346394 500624 346400 500676
rect 346452 500664 346458 500676
rect 349448 500664 349476 500704
rect 351822 500692 351828 500704
rect 351880 500692 351886 500744
rect 354646 500732 354674 501180
rect 354968 501180 365714 501208
rect 354968 500744 354996 501180
rect 371206 500936 371234 501316
rect 416406 500936 416412 500948
rect 365686 500908 367094 500936
rect 371206 500908 416412 500936
rect 365686 500868 365714 500908
rect 364352 500840 365714 500868
rect 367066 500868 367094 500908
rect 416406 500896 416412 500908
rect 416464 500896 416470 500948
rect 416314 500868 416320 500880
rect 367066 500840 416320 500868
rect 364352 500800 364380 500840
rect 416314 500828 416320 500840
rect 416372 500828 416378 500880
rect 416682 500800 416688 500812
rect 364076 500772 364380 500800
rect 364536 500772 416688 500800
rect 364076 500744 364104 500772
rect 354858 500732 354864 500744
rect 354646 500704 354864 500732
rect 354858 500692 354864 500704
rect 354916 500692 354922 500744
rect 354950 500692 354956 500744
rect 355008 500692 355014 500744
rect 364058 500692 364064 500744
rect 364116 500692 364122 500744
rect 364150 500692 364156 500744
rect 364208 500732 364214 500744
rect 364536 500732 364564 500772
rect 416682 500760 416688 500772
rect 416740 500760 416746 500812
rect 364208 500704 364564 500732
rect 364208 500692 364214 500704
rect 364610 500692 364616 500744
rect 364668 500732 364674 500744
rect 416222 500732 416228 500744
rect 364668 500704 416228 500732
rect 364668 500692 364674 500704
rect 416222 500692 416228 500704
rect 416280 500692 416286 500744
rect 416498 500664 416504 500676
rect 346452 500636 349476 500664
rect 349540 500636 416504 500664
rect 346452 500624 346458 500636
rect 196526 500556 196532 500608
rect 196584 500596 196590 500608
rect 203058 500596 203064 500608
rect 196584 500568 203064 500596
rect 196584 500556 196590 500568
rect 203058 500556 203064 500568
rect 203116 500556 203122 500608
rect 203150 500556 203156 500608
rect 203208 500596 203214 500608
rect 238754 500596 238760 500608
rect 203208 500568 238760 500596
rect 203208 500556 203214 500568
rect 238754 500556 238760 500568
rect 238812 500556 238818 500608
rect 343634 500556 343640 500608
rect 343692 500596 343698 500608
rect 349540 500596 349568 500636
rect 416498 500624 416504 500636
rect 416556 500624 416562 500676
rect 343692 500568 349568 500596
rect 343692 500556 343698 500568
rect 349614 500556 349620 500608
rect 349672 500596 349678 500608
rect 416590 500596 416596 500608
rect 349672 500568 416596 500596
rect 349672 500556 349678 500568
rect 416590 500556 416596 500568
rect 416648 500556 416654 500608
rect 174538 500488 174544 500540
rect 174596 500528 174602 500540
rect 219434 500528 219440 500540
rect 174596 500500 219440 500528
rect 174596 500488 174602 500500
rect 219434 500488 219440 500500
rect 219492 500488 219498 500540
rect 336734 500488 336740 500540
rect 336792 500528 336798 500540
rect 418890 500528 418896 500540
rect 336792 500500 418896 500528
rect 336792 500488 336798 500500
rect 418890 500488 418896 500500
rect 418948 500488 418954 500540
rect 196710 500420 196716 500472
rect 196768 500460 196774 500472
rect 203150 500460 203156 500472
rect 196768 500432 203156 500460
rect 196768 500420 196774 500432
rect 203150 500420 203156 500432
rect 203208 500420 203214 500472
rect 203334 500420 203340 500472
rect 203392 500460 203398 500472
rect 242894 500460 242900 500472
rect 203392 500432 242900 500460
rect 203392 500420 203398 500432
rect 242894 500420 242900 500432
rect 242952 500420 242958 500472
rect 333974 500420 333980 500472
rect 334032 500460 334038 500472
rect 419258 500460 419264 500472
rect 334032 500432 419264 500460
rect 334032 500420 334038 500432
rect 419258 500420 419264 500432
rect 419316 500420 419322 500472
rect 195054 500352 195060 500404
rect 195112 500392 195118 500404
rect 241514 500392 241520 500404
rect 195112 500364 241520 500392
rect 195112 500352 195118 500364
rect 241514 500352 241520 500364
rect 241572 500352 241578 500404
rect 329834 500352 329840 500404
rect 329892 500392 329898 500404
rect 419074 500392 419080 500404
rect 329892 500364 419080 500392
rect 329892 500352 329898 500364
rect 419074 500352 419080 500364
rect 419132 500352 419138 500404
rect 196802 500284 196808 500336
rect 196860 500324 196866 500336
rect 244274 500324 244280 500336
rect 196860 500296 244280 500324
rect 196860 500284 196866 500296
rect 244274 500284 244280 500296
rect 244332 500284 244338 500336
rect 327074 500284 327080 500336
rect 327132 500324 327138 500336
rect 418982 500324 418988 500336
rect 327132 500296 418988 500324
rect 327132 500284 327138 500296
rect 418982 500284 418988 500296
rect 419040 500284 419046 500336
rect 196618 500216 196624 500268
rect 196676 500256 196682 500268
rect 254210 500256 254216 500268
rect 196676 500228 202920 500256
rect 196676 500216 196682 500228
rect 202892 500120 202920 500228
rect 206756 500228 254216 500256
rect 206756 500120 206784 500228
rect 254210 500216 254216 500228
rect 254268 500216 254274 500268
rect 324590 500216 324596 500268
rect 324648 500256 324654 500268
rect 418706 500256 418712 500268
rect 324648 500228 418712 500256
rect 324648 500216 324654 500228
rect 418706 500216 418712 500228
rect 418764 500216 418770 500268
rect 213362 500148 213368 500200
rect 213420 500188 213426 500200
rect 215478 500188 215484 500200
rect 213420 500160 215484 500188
rect 213420 500148 213426 500160
rect 215478 500148 215484 500160
rect 215536 500148 215542 500200
rect 340874 500148 340880 500200
rect 340932 500188 340938 500200
rect 349614 500188 349620 500200
rect 340932 500160 349620 500188
rect 340932 500148 340938 500160
rect 349614 500148 349620 500160
rect 349672 500148 349678 500200
rect 351822 500148 351828 500200
rect 351880 500188 351886 500200
rect 357342 500188 357348 500200
rect 351880 500160 357348 500188
rect 351880 500148 351886 500160
rect 357342 500148 357348 500160
rect 357400 500148 357406 500200
rect 357434 500148 357440 500200
rect 357492 500188 357498 500200
rect 415946 500188 415952 500200
rect 357492 500160 415952 500188
rect 357492 500148 357498 500160
rect 415946 500148 415952 500160
rect 416004 500148 416010 500200
rect 202892 500092 206784 500120
rect 207566 500080 207572 500132
rect 207624 500120 207630 500132
rect 215662 500120 215668 500132
rect 207624 500092 215668 500120
rect 207624 500080 207630 500092
rect 215662 500080 215668 500092
rect 215720 500080 215726 500132
rect 351914 500080 351920 500132
rect 351972 500120 351978 500132
rect 364058 500120 364064 500132
rect 351972 500092 364064 500120
rect 351972 500080 351978 500092
rect 364058 500080 364064 500092
rect 364116 500080 364122 500132
rect 357342 500012 357348 500064
rect 357400 500052 357406 500064
rect 364610 500052 364616 500064
rect 357400 500024 364616 500052
rect 357400 500012 357406 500024
rect 364610 500012 364616 500024
rect 364668 500012 364674 500064
rect 19702 499944 19708 499996
rect 19760 499984 19766 499996
rect 20622 499984 20628 499996
rect 19760 499956 20628 499984
rect 19760 499944 19766 499956
rect 20622 499944 20628 499956
rect 20680 499944 20686 499996
rect 15654 499604 15660 499656
rect 15712 499644 15718 499656
rect 17954 499644 17960 499656
rect 15712 499616 17960 499644
rect 15712 499604 15718 499616
rect 17954 499604 17960 499616
rect 18012 499604 18018 499656
rect 15562 499536 15568 499588
rect 15620 499576 15626 499588
rect 19702 499576 19708 499588
rect 15620 499548 19708 499576
rect 15620 499536 15626 499548
rect 19702 499536 19708 499548
rect 19760 499536 19766 499588
rect 17954 499468 17960 499520
rect 18012 499508 18018 499520
rect 18598 499508 18604 499520
rect 18012 499480 18604 499508
rect 18012 499468 18018 499480
rect 18598 499468 18604 499480
rect 18656 499468 18662 499520
rect 244918 499468 244924 499520
rect 244976 499508 244982 499520
rect 389910 499508 389916 499520
rect 244976 499480 389916 499508
rect 244976 499468 244982 499480
rect 389910 499468 389916 499480
rect 389968 499468 389974 499520
rect 20622 499128 20628 499180
rect 20680 499168 20686 499180
rect 51442 499168 51448 499180
rect 20680 499140 51448 499168
rect 20680 499128 20686 499140
rect 51442 499128 51448 499140
rect 51500 499128 51506 499180
rect 18598 499060 18604 499112
rect 18656 499100 18662 499112
rect 53834 499100 53840 499112
rect 18656 499072 53840 499100
rect 18656 499060 18662 499072
rect 53834 499060 53840 499072
rect 53892 499060 53898 499112
rect 194410 499060 194416 499112
rect 194468 499100 194474 499112
rect 249794 499100 249800 499112
rect 194468 499072 249800 499100
rect 194468 499060 194474 499072
rect 249794 499060 249800 499072
rect 249852 499060 249858 499112
rect 17126 498992 17132 499044
rect 17184 499032 17190 499044
rect 60734 499032 60740 499044
rect 17184 499004 60740 499032
rect 17184 498992 17190 499004
rect 60734 498992 60740 499004
rect 60792 498992 60798 499044
rect 193030 498992 193036 499044
rect 193088 499032 193094 499044
rect 251174 499032 251180 499044
rect 193088 499004 251180 499032
rect 193088 498992 193094 499004
rect 251174 498992 251180 499004
rect 251232 498992 251238 499044
rect 7558 498924 7564 498976
rect 7616 498964 7622 498976
rect 219526 498964 219532 498976
rect 7616 498936 219532 498964
rect 7616 498924 7622 498936
rect 219526 498924 219532 498936
rect 219584 498924 219590 498976
rect 261018 498924 261024 498976
rect 261076 498964 261082 498976
rect 381262 498964 381268 498976
rect 261076 498936 381268 498964
rect 261076 498924 261082 498936
rect 381262 498924 381268 498936
rect 381320 498924 381326 498976
rect 17034 498856 17040 498908
rect 17092 498896 17098 498908
rect 59538 498896 59544 498908
rect 17092 498868 59544 498896
rect 17092 498856 17098 498868
rect 59538 498856 59544 498868
rect 59596 498856 59602 498908
rect 207014 498856 207020 498908
rect 207072 498896 207078 498908
rect 558178 498896 558184 498908
rect 207072 498868 558184 498896
rect 207072 498856 207078 498868
rect 558178 498856 558184 498868
rect 558236 498856 558242 498908
rect 19242 498788 19248 498840
rect 19300 498828 19306 498840
rect 385770 498828 385776 498840
rect 19300 498800 385776 498828
rect 19300 498788 19306 498800
rect 385770 498788 385776 498800
rect 385828 498788 385834 498840
rect 419718 498788 419724 498840
rect 419776 498828 419782 498840
rect 454586 498828 454592 498840
rect 419776 498800 454592 498828
rect 419776 498788 419782 498800
rect 454586 498788 454592 498800
rect 454644 498788 454650 498840
rect 15010 498448 15016 498500
rect 15068 498488 15074 498500
rect 34514 498488 34520 498500
rect 15068 498460 34520 498488
rect 15068 498448 15074 498460
rect 34514 498448 34520 498460
rect 34572 498448 34578 498500
rect 16114 498380 16120 498432
rect 16172 498420 16178 498432
rect 44818 498420 44824 498432
rect 16172 498392 44824 498420
rect 16172 498380 16178 498392
rect 44818 498380 44824 498392
rect 44876 498420 44882 498432
rect 45370 498420 45376 498432
rect 44876 498392 45376 498420
rect 44876 498380 44882 498392
rect 45370 498380 45376 498392
rect 45428 498380 45434 498432
rect 16022 498312 16028 498364
rect 16080 498352 16086 498364
rect 18322 498352 18328 498364
rect 16080 498324 18328 498352
rect 16080 498312 16086 498324
rect 18322 498312 18328 498324
rect 18380 498352 18386 498364
rect 58158 498352 58164 498364
rect 18380 498324 58164 498352
rect 18380 498312 18386 498324
rect 58158 498312 58164 498324
rect 58216 498312 58222 498364
rect 15838 498244 15844 498296
rect 15896 498284 15902 498296
rect 55858 498284 55864 498296
rect 15896 498256 55864 498284
rect 15896 498244 15902 498256
rect 55858 498244 55864 498256
rect 55916 498284 55922 498296
rect 57882 498284 57888 498296
rect 55916 498256 57888 498284
rect 55916 498244 55922 498256
rect 57882 498244 57888 498256
rect 57940 498244 57946 498296
rect 14826 498176 14832 498228
rect 14884 498216 14890 498228
rect 15010 498216 15016 498228
rect 14884 498188 15016 498216
rect 14884 498176 14890 498188
rect 15010 498176 15016 498188
rect 15068 498176 15074 498228
rect 16298 498176 16304 498228
rect 16356 498216 16362 498228
rect 57054 498216 57060 498228
rect 16356 498188 57060 498216
rect 16356 498176 16362 498188
rect 57054 498176 57060 498188
rect 57112 498176 57118 498228
rect 389358 498176 389364 498228
rect 389416 498216 389422 498228
rect 389910 498216 389916 498228
rect 389416 498188 389916 498216
rect 389416 498176 389422 498188
rect 389910 498176 389916 498188
rect 389968 498176 389974 498228
rect 19058 498108 19064 498160
rect 19116 498148 19122 498160
rect 52178 498148 52184 498160
rect 19116 498120 52184 498148
rect 19116 498108 19122 498120
rect 52178 498108 52184 498120
rect 52236 498108 52242 498160
rect 59538 498108 59544 498160
rect 59596 498148 59602 498160
rect 78122 498148 78128 498160
rect 59596 498120 78128 498148
rect 59596 498108 59602 498120
rect 78122 498108 78128 498120
rect 78180 498108 78186 498160
rect 196434 498108 196440 498160
rect 196492 498148 196498 498160
rect 228542 498148 228548 498160
rect 196492 498120 228548 498148
rect 196492 498108 196498 498120
rect 228542 498108 228548 498120
rect 228600 498108 228606 498160
rect 302234 498108 302240 498160
rect 302292 498148 302298 498160
rect 413278 498148 413284 498160
rect 302292 498120 413284 498148
rect 302292 498108 302298 498120
rect 413278 498108 413284 498120
rect 413336 498108 413342 498160
rect 454586 498108 454592 498160
rect 454644 498148 454650 498160
rect 473354 498148 473360 498160
rect 454644 498120 473360 498148
rect 454644 498108 454650 498120
rect 473354 498108 473360 498120
rect 473412 498108 473418 498160
rect 16390 498040 16396 498092
rect 16448 498080 16454 498092
rect 46842 498080 46848 498092
rect 16448 498052 46848 498080
rect 16448 498040 16454 498052
rect 46842 498040 46848 498052
rect 46900 498040 46906 498092
rect 195514 498040 195520 498092
rect 195572 498080 195578 498092
rect 228634 498080 228640 498092
rect 195572 498052 228640 498080
rect 195572 498040 195578 498052
rect 228634 498040 228640 498052
rect 228692 498040 228698 498092
rect 259638 498040 259644 498092
rect 259696 498080 259702 498092
rect 378502 498080 378508 498092
rect 259696 498052 378508 498080
rect 259696 498040 259702 498052
rect 378502 498040 378508 498052
rect 378560 498040 378566 498092
rect 19978 497972 19984 498024
rect 20036 498012 20042 498024
rect 48682 498012 48688 498024
rect 20036 497984 48688 498012
rect 20036 497972 20042 497984
rect 48682 497972 48688 497984
rect 48740 498012 48746 498024
rect 49602 498012 49608 498024
rect 48740 497984 49608 498012
rect 48740 497972 48746 497984
rect 49602 497972 49608 497984
rect 49660 497972 49666 498024
rect 195238 497972 195244 498024
rect 195296 498012 195302 498024
rect 238846 498012 238852 498024
rect 195296 497984 238852 498012
rect 195296 497972 195302 497984
rect 238846 497972 238852 497984
rect 238904 497972 238910 498024
rect 258166 497972 258172 498024
rect 258224 498012 258230 498024
rect 377674 498012 377680 498024
rect 258224 497984 377680 498012
rect 258224 497972 258230 497984
rect 377674 497972 377680 497984
rect 377732 497972 377738 498024
rect 18414 497904 18420 497956
rect 18472 497944 18478 497956
rect 39666 497944 39672 497956
rect 18472 497916 39672 497944
rect 18472 497904 18478 497916
rect 39666 497904 39672 497916
rect 39724 497904 39730 497956
rect 52454 497904 52460 497956
rect 52512 497944 52518 497956
rect 53466 497944 53472 497956
rect 52512 497916 53472 497944
rect 52512 497904 52518 497916
rect 53466 497904 53472 497916
rect 53524 497944 53530 497956
rect 71958 497944 71964 497956
rect 53524 497916 71964 497944
rect 53524 497904 53530 497916
rect 71958 497904 71964 497916
rect 72016 497904 72022 497956
rect 199194 497904 199200 497956
rect 199252 497944 199258 497956
rect 259454 497944 259460 497956
rect 199252 497916 259460 497944
rect 199252 497904 199258 497916
rect 259454 497904 259460 497916
rect 259512 497904 259518 497956
rect 259546 497904 259552 497956
rect 259604 497944 259610 497956
rect 379790 497944 379796 497956
rect 259604 497916 379796 497944
rect 259604 497904 259610 497916
rect 379790 497904 379796 497916
rect 379848 497904 379854 497956
rect 34514 497836 34520 497888
rect 34572 497876 34578 497888
rect 47578 497876 47584 497888
rect 34572 497848 47584 497876
rect 34572 497836 34578 497848
rect 47578 497836 47584 497848
rect 47636 497876 47642 497888
rect 48222 497876 48228 497888
rect 47636 497848 48228 497876
rect 47636 497836 47642 497848
rect 48222 497836 48228 497848
rect 48280 497836 48286 497888
rect 51442 497836 51448 497888
rect 51500 497876 51506 497888
rect 69658 497876 69664 497888
rect 51500 497848 69664 497876
rect 51500 497836 51506 497848
rect 69658 497836 69664 497848
rect 69716 497836 69722 497888
rect 197078 497836 197084 497888
rect 197136 497876 197142 497888
rect 256694 497876 256700 497888
rect 197136 497848 256700 497876
rect 197136 497836 197142 497848
rect 256694 497836 256700 497848
rect 256752 497836 256758 497888
rect 258258 497836 258264 497888
rect 258316 497876 258322 497888
rect 379606 497876 379612 497888
rect 258316 497848 379612 497876
rect 258316 497836 258322 497848
rect 379606 497836 379612 497848
rect 379664 497836 379670 497888
rect 19886 497768 19892 497820
rect 19944 497808 19950 497820
rect 37182 497808 37188 497820
rect 19944 497780 37188 497808
rect 19944 497768 19950 497780
rect 37182 497768 37188 497780
rect 37240 497808 37246 497820
rect 42794 497808 42800 497820
rect 37240 497780 42800 497808
rect 37240 497768 37246 497780
rect 42794 497768 42800 497780
rect 42852 497768 42858 497820
rect 57882 497768 57888 497820
rect 57940 497808 57946 497820
rect 73982 497808 73988 497820
rect 57940 497780 73988 497808
rect 57940 497768 57946 497780
rect 73982 497768 73988 497780
rect 74040 497768 74046 497820
rect 195146 497768 195152 497820
rect 195204 497808 195210 497820
rect 255406 497808 255412 497820
rect 195204 497780 255412 497808
rect 195204 497768 195210 497780
rect 255406 497768 255412 497780
rect 255464 497768 255470 497820
rect 256786 497768 256792 497820
rect 256844 497808 256850 497820
rect 378410 497808 378416 497820
rect 256844 497780 378416 497808
rect 256844 497768 256850 497780
rect 378410 497768 378416 497780
rect 378468 497768 378474 497820
rect 19150 497700 19156 497752
rect 19208 497740 19214 497752
rect 36170 497740 36176 497752
rect 19208 497712 36176 497740
rect 19208 497700 19214 497712
rect 36170 497700 36176 497712
rect 36228 497740 36234 497752
rect 38654 497740 38660 497752
rect 36228 497712 38660 497740
rect 36228 497700 36234 497712
rect 38654 497700 38660 497712
rect 38712 497700 38718 497752
rect 53834 497700 53840 497752
rect 53892 497740 53898 497752
rect 73154 497740 73160 497752
rect 53892 497712 73160 497740
rect 53892 497700 53898 497712
rect 73154 497700 73160 497712
rect 73212 497700 73218 497752
rect 201218 497700 201224 497752
rect 201276 497740 201282 497752
rect 247126 497740 247132 497752
rect 201276 497712 247132 497740
rect 201276 497700 201282 497712
rect 247126 497700 247132 497712
rect 247184 497700 247190 497752
rect 255590 497700 255596 497752
rect 255648 497740 255654 497752
rect 378318 497740 378324 497752
rect 255648 497712 378324 497740
rect 255648 497700 255654 497712
rect 378318 497700 378324 497712
rect 378376 497700 378382 497752
rect 445294 497700 445300 497752
rect 445352 497740 445358 497752
rect 463694 497740 463700 497752
rect 445352 497712 463700 497740
rect 445352 497700 445358 497712
rect 463694 497700 463700 497712
rect 463752 497700 463758 497752
rect 60642 497632 60648 497684
rect 60700 497672 60706 497684
rect 79410 497672 79416 497684
rect 60700 497644 79416 497672
rect 60700 497632 60706 497644
rect 79410 497632 79416 497644
rect 79468 497632 79474 497684
rect 196986 497632 196992 497684
rect 197044 497672 197050 497684
rect 244366 497672 244372 497684
rect 197044 497644 244372 497672
rect 197044 497632 197050 497644
rect 244366 497632 244372 497644
rect 244424 497632 244430 497684
rect 254026 497632 254032 497684
rect 254084 497672 254090 497684
rect 378226 497672 378232 497684
rect 254084 497644 378232 497672
rect 254084 497632 254090 497644
rect 378226 497632 378232 497644
rect 378284 497632 378290 497684
rect 419902 497632 419908 497684
rect 419960 497672 419966 497684
rect 437474 497672 437480 497684
rect 419960 497644 437480 497672
rect 419960 497632 419966 497644
rect 437474 497632 437480 497644
rect 437532 497632 437538 497684
rect 444190 497632 444196 497684
rect 444248 497672 444254 497684
rect 462314 497672 462320 497684
rect 444248 497644 462320 497672
rect 444248 497632 444254 497644
rect 462314 497632 462320 497644
rect 462372 497632 462378 497684
rect 462498 497632 462504 497684
rect 462556 497672 462562 497684
rect 476114 497672 476120 497684
rect 462556 497644 476120 497672
rect 462556 497632 462562 497644
rect 476114 497632 476120 497644
rect 476172 497632 476178 497684
rect 16022 497564 16028 497616
rect 16080 497604 16086 497616
rect 19978 497604 19984 497616
rect 16080 497576 19984 497604
rect 16080 497564 16086 497576
rect 19978 497564 19984 497576
rect 20036 497564 20042 497616
rect 22094 497564 22100 497616
rect 22152 497604 22158 497616
rect 40586 497604 40592 497616
rect 22152 497576 40592 497604
rect 22152 497564 22158 497576
rect 40586 497564 40592 497576
rect 40644 497564 40650 497616
rect 44818 497564 44824 497616
rect 44876 497604 44882 497616
rect 64138 497604 64144 497616
rect 44876 497576 64144 497604
rect 44876 497564 44882 497576
rect 64138 497564 64144 497576
rect 64196 497564 64202 497616
rect 196894 497564 196900 497616
rect 196952 497604 196958 497616
rect 241606 497604 241612 497616
rect 196952 497576 241612 497604
rect 196952 497564 196958 497576
rect 241606 497564 241612 497576
rect 241664 497564 241670 497616
rect 242986 497564 242992 497616
rect 243044 497604 243050 497616
rect 381170 497604 381176 497616
rect 243044 497576 381176 497604
rect 243044 497564 243050 497576
rect 381170 497564 381176 497576
rect 381228 497564 381234 497616
rect 419810 497564 419816 497616
rect 419868 497604 419874 497616
rect 438854 497604 438860 497616
rect 419868 497576 438860 497604
rect 419868 497564 419874 497576
rect 438854 497564 438860 497576
rect 438912 497564 438918 497616
rect 462038 497564 462044 497616
rect 462096 497604 462102 497616
rect 474734 497604 474740 497616
rect 462096 497576 474740 497604
rect 462096 497564 462102 497576
rect 474734 497564 474740 497576
rect 474792 497564 474798 497616
rect 19794 497496 19800 497548
rect 19852 497536 19858 497548
rect 43438 497536 43444 497548
rect 19852 497508 43444 497536
rect 19852 497496 19858 497508
rect 43438 497496 43444 497508
rect 43496 497496 43502 497548
rect 49602 497496 49608 497548
rect 49660 497536 49666 497548
rect 67634 497536 67640 497548
rect 49660 497508 67640 497536
rect 49660 497496 49666 497508
rect 67634 497496 67640 497508
rect 67692 497536 67698 497548
rect 68922 497536 68928 497548
rect 67692 497508 68928 497536
rect 67692 497496 67698 497508
rect 68922 497496 68928 497508
rect 68980 497496 68986 497548
rect 195330 497496 195336 497548
rect 195388 497536 195394 497548
rect 240134 497536 240140 497548
rect 195388 497508 240140 497536
rect 195388 497496 195394 497508
rect 240134 497496 240140 497508
rect 240192 497496 240198 497548
rect 240226 497496 240232 497548
rect 240284 497536 240290 497548
rect 379698 497536 379704 497548
rect 240284 497508 379704 497536
rect 240284 497496 240290 497508
rect 379698 497496 379704 497508
rect 379756 497496 379762 497548
rect 417970 497496 417976 497548
rect 418028 497536 418034 497548
rect 451274 497536 451280 497548
rect 418028 497508 451280 497536
rect 418028 497496 418034 497508
rect 451274 497496 451280 497508
rect 451332 497536 451338 497548
rect 469214 497536 469220 497548
rect 451332 497508 469220 497536
rect 451332 497496 451338 497508
rect 469214 497496 469220 497508
rect 469272 497496 469278 497548
rect 15010 497428 15016 497480
rect 15068 497468 15074 497480
rect 52454 497468 52460 497480
rect 15068 497440 52460 497468
rect 15068 497428 15074 497440
rect 52454 497428 52460 497440
rect 52512 497428 52518 497480
rect 70394 497428 70400 497480
rect 70452 497468 70458 497480
rect 71222 497468 71228 497480
rect 70452 497440 71228 497468
rect 70452 497428 70458 497440
rect 71222 497428 71228 497440
rect 71280 497468 71286 497480
rect 313274 497468 313280 497480
rect 71280 497440 313280 497468
rect 71280 497428 71286 497440
rect 313274 497428 313280 497440
rect 313332 497428 313338 497480
rect 334894 497428 334900 497480
rect 334952 497468 334958 497480
rect 391934 497468 391940 497480
rect 334952 497440 391940 497468
rect 334952 497428 334958 497440
rect 391934 497428 391940 497440
rect 391992 497428 391998 497480
rect 418062 497428 418068 497480
rect 418120 497468 418126 497480
rect 452378 497468 452384 497480
rect 418120 497440 452384 497468
rect 418120 497428 418126 497440
rect 452378 497428 452384 497440
rect 452436 497468 452442 497480
rect 470870 497468 470876 497480
rect 452436 497440 470876 497468
rect 452436 497428 452442 497440
rect 470870 497428 470876 497440
rect 470928 497428 470934 497480
rect 197170 497360 197176 497412
rect 197228 497400 197234 497412
rect 228726 497400 228732 497412
rect 197228 497372 228732 497400
rect 197228 497360 197234 497372
rect 228726 497360 228732 497372
rect 228784 497360 228790 497412
rect 360470 497360 360476 497412
rect 360528 497400 360534 497412
rect 416130 497400 416136 497412
rect 360528 497372 416136 497400
rect 360528 497360 360534 497372
rect 416130 497360 416136 497372
rect 416188 497360 416194 497412
rect 449158 497360 449164 497412
rect 449216 497400 449222 497412
rect 466454 497400 466460 497412
rect 449216 497372 466460 497400
rect 449216 497360 449222 497372
rect 466454 497360 466460 497372
rect 466512 497360 466518 497412
rect 450538 497292 450544 497344
rect 450596 497332 450602 497344
rect 467834 497332 467840 497344
rect 450596 497304 467840 497332
rect 450596 497292 450602 497304
rect 467834 497292 467840 497304
rect 467892 497292 467898 497344
rect 447778 497224 447784 497276
rect 447836 497264 447842 497276
rect 465074 497264 465080 497276
rect 447836 497236 465080 497264
rect 447836 497224 447842 497236
rect 465074 497224 465080 497236
rect 465132 497224 465138 497276
rect 20622 497156 20628 497208
rect 20680 497196 20686 497208
rect 44174 497196 44180 497208
rect 20680 497168 44180 497196
rect 20680 497156 20686 497168
rect 44174 497156 44180 497168
rect 44232 497196 44238 497208
rect 62758 497196 62764 497208
rect 44232 497168 62764 497196
rect 44232 497156 44238 497168
rect 62758 497156 62764 497168
rect 62816 497156 62822 497208
rect 443638 497156 443644 497208
rect 443696 497196 443702 497208
rect 461118 497196 461124 497208
rect 443696 497168 461124 497196
rect 443696 497156 443702 497168
rect 461118 497156 461124 497168
rect 461176 497156 461182 497208
rect 43438 497088 43444 497140
rect 43496 497128 43502 497140
rect 61838 497128 61844 497140
rect 43496 497100 61844 497128
rect 43496 497088 43502 497100
rect 61838 497088 61844 497100
rect 61896 497088 61902 497140
rect 78122 497088 78128 497140
rect 78180 497128 78186 497140
rect 79318 497128 79324 497140
rect 78180 497100 79324 497128
rect 78180 497088 78186 497100
rect 79318 497088 79324 497100
rect 79376 497088 79382 497140
rect 456058 497088 456064 497140
rect 456116 497128 456122 497140
rect 473354 497128 473360 497140
rect 456116 497100 473360 497128
rect 456116 497088 456122 497100
rect 473354 497088 473360 497100
rect 473412 497088 473418 497140
rect 50246 497060 50252 497072
rect 45526 497032 50252 497060
rect 45526 496992 45554 497032
rect 50246 497020 50252 497032
rect 50304 497060 50310 497072
rect 68278 497060 68284 497072
rect 50304 497032 68284 497060
rect 50304 497020 50310 497032
rect 68278 497020 68284 497032
rect 68336 497020 68342 497072
rect 71958 497020 71964 497072
rect 72016 497060 72022 497072
rect 319438 497060 319444 497072
rect 72016 497032 319444 497060
rect 72016 497020 72022 497032
rect 319438 497020 319444 497032
rect 319496 497020 319502 497072
rect 446674 497020 446680 497072
rect 446732 497060 446738 497072
rect 465074 497060 465080 497072
rect 446732 497032 465080 497060
rect 446732 497020 446738 497032
rect 465074 497020 465080 497032
rect 465132 497020 465138 497072
rect 35866 496964 45554 496992
rect 16482 496748 16488 496800
rect 16540 496788 16546 496800
rect 34514 496788 34520 496800
rect 16540 496760 34520 496788
rect 16540 496748 16546 496760
rect 34514 496748 34520 496760
rect 34572 496788 34578 496800
rect 35866 496788 35894 496964
rect 52178 496952 52184 497004
rect 52236 496992 52242 497004
rect 52454 496992 52460 497004
rect 52236 496964 52460 496992
rect 52236 496952 52242 496964
rect 52454 496952 52460 496964
rect 52512 496992 52518 497004
rect 70394 496992 70400 497004
rect 52512 496964 70400 496992
rect 52512 496952 52518 496964
rect 70394 496952 70400 496964
rect 70452 496952 70458 497004
rect 313274 496952 313280 497004
rect 313332 496992 313338 497004
rect 315298 496992 315304 497004
rect 313332 496964 315304 496992
rect 313332 496952 313338 496964
rect 315298 496952 315304 496964
rect 315356 496992 315362 497004
rect 315356 496964 417372 496992
rect 315356 496952 315362 496964
rect 417344 496936 417372 496964
rect 459554 496952 459560 497004
rect 459612 496992 459618 497004
rect 460566 496992 460572 497004
rect 459612 496964 460572 496992
rect 459612 496952 459618 496964
rect 460566 496952 460572 496964
rect 460624 496992 460630 497004
rect 478874 496992 478880 497004
rect 460624 496964 478880 496992
rect 460624 496952 460630 496964
rect 478874 496952 478880 496964
rect 478932 496952 478938 497004
rect 39666 496884 39672 496936
rect 39724 496924 39730 496936
rect 44174 496924 44180 496936
rect 39724 496896 44180 496924
rect 39724 496884 39730 496896
rect 44174 496884 44180 496896
rect 44232 496884 44238 496936
rect 48222 496884 48228 496936
rect 48280 496924 48286 496936
rect 66254 496924 66260 496936
rect 48280 496896 66260 496924
rect 48280 496884 48286 496896
rect 66254 496884 66260 496896
rect 66312 496924 66318 496936
rect 66898 496924 66904 496936
rect 66312 496896 66904 496924
rect 66312 496884 66318 496896
rect 66898 496884 66904 496896
rect 66956 496884 66962 496936
rect 68922 496884 68928 496936
rect 68980 496924 68986 496936
rect 301498 496924 301504 496936
rect 68980 496896 301504 496924
rect 68980 496884 68986 496896
rect 301498 496884 301504 496896
rect 301556 496884 301562 496936
rect 311158 496884 311164 496936
rect 311216 496924 311222 496936
rect 311216 496896 412634 496924
rect 311216 496884 311222 496896
rect 40586 496816 40592 496868
rect 40644 496856 40650 496868
rect 43438 496856 43444 496868
rect 40644 496828 43444 496856
rect 40644 496816 40650 496828
rect 43438 496816 43444 496828
rect 43496 496816 43502 496868
rect 46842 496816 46848 496868
rect 46900 496856 46906 496868
rect 65518 496856 65524 496868
rect 46900 496828 65524 496856
rect 46900 496816 46906 496828
rect 65518 496816 65524 496828
rect 65576 496816 65582 496868
rect 412606 496856 412634 496896
rect 417326 496884 417332 496936
rect 417384 496924 417390 496936
rect 418062 496924 418068 496936
rect 417384 496896 418068 496924
rect 417384 496884 417390 496896
rect 418062 496884 418068 496896
rect 418120 496884 418126 496936
rect 453298 496884 453304 496936
rect 453356 496924 453362 496936
rect 471974 496924 471980 496936
rect 453356 496896 471980 496924
rect 453356 496884 453362 496896
rect 471974 496884 471980 496896
rect 472032 496884 472038 496936
rect 417234 496856 417240 496868
rect 412606 496828 417240 496856
rect 417234 496816 417240 496828
rect 417292 496856 417298 496868
rect 417970 496856 417976 496868
rect 417292 496828 417976 496856
rect 417292 496816 417298 496828
rect 417970 496816 417976 496828
rect 418028 496816 418034 496868
rect 420730 496816 420736 496868
rect 420788 496856 420794 496868
rect 436094 496856 436100 496868
rect 420788 496828 436100 496856
rect 420788 496816 420794 496828
rect 436094 496816 436100 496828
rect 436152 496816 436158 496868
rect 458818 496816 458824 496868
rect 458876 496856 458882 496868
rect 459462 496856 459468 496868
rect 458876 496828 459468 496856
rect 458876 496816 458882 496828
rect 459462 496816 459468 496828
rect 459520 496856 459526 496868
rect 477494 496856 477500 496868
rect 459520 496828 477500 496856
rect 459520 496816 459526 496828
rect 477494 496816 477500 496828
rect 477552 496816 477558 496868
rect 34572 496760 35894 496788
rect 34572 496748 34578 496760
rect 419994 496748 420000 496800
rect 420052 496788 420058 496800
rect 459554 496788 459560 496800
rect 420052 496760 459560 496788
rect 420052 496748 420058 496760
rect 459554 496748 459560 496760
rect 459612 496748 459618 496800
rect 15102 496680 15108 496732
rect 15160 496720 15166 496732
rect 19794 496720 19800 496732
rect 15160 496692 19800 496720
rect 15160 496680 15166 496692
rect 19794 496680 19800 496692
rect 19852 496720 19858 496732
rect 20622 496720 20628 496732
rect 19852 496692 20628 496720
rect 19852 496680 19858 496692
rect 20622 496680 20628 496692
rect 20680 496680 20686 496732
rect 419442 496680 419448 496732
rect 419500 496720 419506 496732
rect 445754 496720 445760 496732
rect 419500 496692 445760 496720
rect 419500 496680 419506 496692
rect 445754 496680 445760 496692
rect 445812 496720 445818 496732
rect 446674 496720 446680 496732
rect 445812 496692 446680 496720
rect 445812 496680 445818 496692
rect 446674 496680 446680 496692
rect 446732 496680 446738 496732
rect 201586 496204 201592 496256
rect 201644 496244 201650 496256
rect 235258 496244 235264 496256
rect 201644 496216 235264 496244
rect 201644 496204 201650 496216
rect 235258 496204 235264 496216
rect 235316 496204 235322 496256
rect 212718 496136 212724 496188
rect 212776 496176 212782 496188
rect 389818 496176 389824 496188
rect 212776 496148 389824 496176
rect 212776 496136 212782 496148
rect 389818 496136 389824 496148
rect 389876 496136 389882 496188
rect 63678 496068 63684 496120
rect 63736 496108 63742 496120
rect 304994 496108 305000 496120
rect 63736 496080 305000 496108
rect 63736 496068 63742 496080
rect 304994 496068 305000 496080
rect 305052 496068 305058 496120
rect 316034 496068 316040 496120
rect 316092 496108 316098 496120
rect 470778 496108 470784 496120
rect 316092 496080 470784 496108
rect 316092 496068 316098 496080
rect 470778 496068 470784 496080
rect 470836 496068 470842 496120
rect 338758 495524 338764 495576
rect 338816 495564 338822 495576
rect 418154 495564 418160 495576
rect 338816 495536 418160 495564
rect 338816 495524 338822 495536
rect 418154 495524 418160 495536
rect 418212 495564 418218 495576
rect 419994 495564 420000 495576
rect 418212 495536 420000 495564
rect 418212 495524 418218 495536
rect 419994 495524 420000 495536
rect 420052 495524 420058 495576
rect 278038 495456 278044 495508
rect 278096 495496 278102 495508
rect 418706 495496 418712 495508
rect 278096 495468 418712 495496
rect 278096 495456 278102 495468
rect 418706 495456 418712 495468
rect 418764 495456 418770 495508
rect 286318 495184 286324 495236
rect 286376 495224 286382 495236
rect 413738 495224 413744 495236
rect 286376 495196 413744 495224
rect 286376 495184 286382 495196
rect 413738 495184 413744 495196
rect 413796 495224 413802 495236
rect 415302 495224 415308 495236
rect 413796 495196 415308 495224
rect 413796 495184 413802 495196
rect 415302 495184 415308 495196
rect 415360 495184 415366 495236
rect 252830 495116 252836 495168
rect 252888 495156 252894 495168
rect 381078 495156 381084 495168
rect 252888 495128 381084 495156
rect 252888 495116 252894 495128
rect 381078 495116 381084 495128
rect 381136 495116 381142 495168
rect 248414 495048 248420 495100
rect 248472 495088 248478 495100
rect 377582 495088 377588 495100
rect 248472 495060 377588 495088
rect 248472 495048 248478 495060
rect 377582 495048 377588 495060
rect 377640 495048 377646 495100
rect 194502 494980 194508 495032
rect 194560 495020 194566 495032
rect 232498 495020 232504 495032
rect 194560 494992 232504 495020
rect 194560 494980 194566 494992
rect 232498 494980 232504 494992
rect 232556 494980 232562 495032
rect 249886 494980 249892 495032
rect 249944 495020 249950 495032
rect 379514 495020 379520 495032
rect 249944 494992 379520 495020
rect 249944 494980 249950 494992
rect 379514 494980 379520 494992
rect 379572 494980 379578 495032
rect 193122 494912 193128 494964
rect 193180 494952 193186 494964
rect 232590 494952 232596 494964
rect 193180 494924 232596 494952
rect 193180 494912 193186 494924
rect 232590 494912 232596 494924
rect 232648 494912 232654 494964
rect 251266 494912 251272 494964
rect 251324 494952 251330 494964
rect 380986 494952 380992 494964
rect 251324 494924 380992 494952
rect 251324 494912 251330 494924
rect 380986 494912 380992 494924
rect 381044 494912 381050 494964
rect 106090 494844 106096 494896
rect 106148 494884 106154 494896
rect 360286 494884 360292 494896
rect 106148 494856 360292 494884
rect 106148 494844 106154 494856
rect 360286 494844 360292 494856
rect 360344 494844 360350 494896
rect 415302 494844 415308 494896
rect 415360 494884 415366 494896
rect 444190 494884 444196 494896
rect 415360 494856 444196 494884
rect 415360 494844 415366 494856
rect 444190 494844 444196 494856
rect 444248 494844 444254 494896
rect 16942 494776 16948 494828
rect 17000 494816 17006 494828
rect 304350 494816 304356 494828
rect 17000 494788 304356 494816
rect 17000 494776 17006 494788
rect 304350 494776 304356 494788
rect 304408 494776 304414 494828
rect 319070 494776 319076 494828
rect 319128 494816 319134 494828
rect 473538 494816 473544 494828
rect 319128 494788 473544 494816
rect 319128 494776 319134 494788
rect 473538 494776 473544 494788
rect 473596 494776 473602 494828
rect 207106 494708 207112 494760
rect 207164 494748 207170 494760
rect 571978 494748 571984 494760
rect 207164 494720 571984 494748
rect 207164 494708 207170 494720
rect 571978 494708 571984 494720
rect 572036 494708 572042 494760
rect 48314 493484 48320 493536
rect 48372 493524 48378 493536
rect 280246 493524 280252 493536
rect 48372 493496 280252 493524
rect 48372 493484 48378 493496
rect 280246 493484 280252 493496
rect 280304 493484 280310 493536
rect 41874 493416 41880 493468
rect 41932 493456 41938 493468
rect 293954 493456 293960 493468
rect 41932 493428 293960 493456
rect 41932 493416 41938 493428
rect 293954 493416 293960 493428
rect 294012 493416 294018 493468
rect 325970 493416 325976 493468
rect 326028 493456 326034 493468
rect 477586 493456 477592 493468
rect 326028 493428 477592 493456
rect 326028 493416 326034 493428
rect 477586 493416 477592 493428
rect 477644 493416 477650 493468
rect 100938 493348 100944 493400
rect 100996 493388 101002 493400
rect 354766 493388 354772 493400
rect 100996 493360 354772 493388
rect 100996 493348 101002 493360
rect 354766 493348 354772 493360
rect 354824 493348 354830 493400
rect 208394 493280 208400 493332
rect 208452 493320 208458 493332
rect 569218 493320 569224 493332
rect 208452 493292 569224 493320
rect 208452 493280 208458 493292
rect 569218 493280 569224 493292
rect 569276 493280 569282 493332
rect 293954 492668 293960 492720
rect 294012 492708 294018 492720
rect 294230 492708 294236 492720
rect 294012 492680 294236 492708
rect 294012 492668 294018 492680
rect 294230 492668 294236 492680
rect 294288 492708 294294 492720
rect 416682 492708 416688 492720
rect 294288 492680 416688 492708
rect 294288 492668 294294 492680
rect 416682 492668 416688 492680
rect 416740 492668 416746 492720
rect 416774 492600 416780 492652
rect 416832 492640 416838 492652
rect 417786 492640 417792 492652
rect 416832 492612 417792 492640
rect 416832 492600 416838 492612
rect 417786 492600 417792 492612
rect 417844 492640 417850 492652
rect 456886 492640 456892 492652
rect 417844 492612 456892 492640
rect 417844 492600 417850 492612
rect 456886 492600 456892 492612
rect 456944 492600 456950 492652
rect 208486 492056 208492 492108
rect 208544 492096 208550 492108
rect 382918 492096 382924 492108
rect 208544 492068 382924 492096
rect 208544 492056 208550 492068
rect 382918 492056 382924 492068
rect 382976 492056 382982 492108
rect 73706 491988 73712 492040
rect 73764 492028 73770 492040
rect 320266 492028 320272 492040
rect 73764 492000 320272 492028
rect 73764 491988 73770 492000
rect 320266 491988 320272 492000
rect 320324 491988 320330 492040
rect 328454 491988 328460 492040
rect 328512 492028 328518 492040
rect 480530 492028 480536 492040
rect 328512 492000 480536 492028
rect 328512 491988 328518 492000
rect 480530 491988 480536 492000
rect 480588 491988 480594 492040
rect 108850 491920 108856 491972
rect 108908 491960 108914 491972
rect 363230 491960 363236 491972
rect 108908 491932 363236 491960
rect 108908 491920 108914 491932
rect 363230 491920 363236 491932
rect 363288 491920 363294 491972
rect 329098 491308 329104 491360
rect 329156 491348 329162 491360
rect 417786 491348 417792 491360
rect 329156 491320 417792 491348
rect 329156 491308 329162 491320
rect 417786 491308 417792 491320
rect 417844 491308 417850 491360
rect 292482 490832 292488 490884
rect 292540 490872 292546 490884
rect 413830 490872 413836 490884
rect 292540 490844 413836 490872
rect 292540 490832 292546 490844
rect 413830 490832 413836 490844
rect 413888 490872 413894 490884
rect 415210 490872 415216 490884
rect 413888 490844 415216 490872
rect 413888 490832 413894 490844
rect 415210 490832 415216 490844
rect 415268 490832 415274 490884
rect 209774 490764 209780 490816
rect 209832 490804 209838 490816
rect 385678 490804 385684 490816
rect 209832 490776 385684 490804
rect 209832 490764 209838 490776
rect 385678 490764 385684 490776
rect 385736 490764 385742 490816
rect 61838 490696 61844 490748
rect 61896 490736 61902 490748
rect 281810 490736 281816 490748
rect 61896 490708 281816 490736
rect 61896 490696 61902 490708
rect 281810 490696 281816 490708
rect 281868 490696 281874 490748
rect 301038 490696 301044 490748
rect 301096 490736 301102 490748
rect 460934 490736 460940 490748
rect 301096 490708 460940 490736
rect 301096 490696 301102 490708
rect 460934 490696 460940 490708
rect 460992 490696 460998 490748
rect 68554 490628 68560 490680
rect 68612 490668 68618 490680
rect 313274 490668 313280 490680
rect 68612 490640 313280 490668
rect 68612 490628 68618 490640
rect 313274 490628 313280 490640
rect 313332 490628 313338 490680
rect 415210 490628 415216 490680
rect 415268 490668 415274 490680
rect 445294 490668 445300 490680
rect 415268 490640 445300 490668
rect 415268 490628 415274 490640
rect 445294 490628 445300 490640
rect 445352 490628 445358 490680
rect 76834 490560 76840 490612
rect 76892 490600 76898 490612
rect 322934 490600 322940 490612
rect 76892 490572 322940 490600
rect 76892 490560 76898 490572
rect 322934 490560 322940 490572
rect 322992 490560 322998 490612
rect 342254 490560 342260 490612
rect 342312 490600 342318 490612
rect 490466 490600 490472 490612
rect 342312 490572 490472 490600
rect 342312 490560 342318 490572
rect 490466 490560 490472 490572
rect 490524 490560 490530 490612
rect 64138 489812 64144 489864
rect 64196 489852 64202 489864
rect 291194 489852 291200 489864
rect 64196 489824 291200 489852
rect 64196 489812 64202 489824
rect 291194 489812 291200 489824
rect 291252 489812 291258 489864
rect 159450 489268 159456 489320
rect 159508 489308 159514 489320
rect 349246 489308 349252 489320
rect 159508 489280 349252 489308
rect 159508 489268 159514 489280
rect 349246 489268 349252 489280
rect 349304 489268 349310 489320
rect 37274 489200 37280 489252
rect 37332 489240 37338 489252
rect 280798 489240 280804 489252
rect 37332 489212 280804 489240
rect 37332 489200 37338 489212
rect 280798 489200 280804 489212
rect 280856 489200 280862 489252
rect 287054 489200 287060 489252
rect 287112 489240 287118 489252
rect 452654 489240 452660 489252
rect 287112 489212 452660 489240
rect 287112 489200 287118 489212
rect 452654 489200 452660 489212
rect 452712 489200 452718 489252
rect 78582 489132 78588 489184
rect 78640 489172 78646 489184
rect 325786 489172 325792 489184
rect 78640 489144 325792 489172
rect 78640 489132 78646 489144
rect 325786 489132 325792 489144
rect 325844 489132 325850 489184
rect 353294 489132 353300 489184
rect 353352 489172 353358 489184
rect 500954 489172 500960 489184
rect 353352 489144 500960 489172
rect 353352 489132 353358 489144
rect 500954 489132 500960 489144
rect 501012 489132 501018 489184
rect 291194 488724 291200 488776
rect 291252 488764 291258 488776
rect 292482 488764 292488 488776
rect 291252 488736 292488 488764
rect 291252 488724 291258 488736
rect 292482 488724 292488 488736
rect 292540 488724 292546 488776
rect 417878 488452 417884 488504
rect 417936 488492 417942 488504
rect 456058 488492 456064 488504
rect 417936 488464 456064 488492
rect 417936 488452 417942 488464
rect 456058 488452 456064 488464
rect 456116 488452 456122 488504
rect 292850 487976 292856 488028
rect 292908 488016 292914 488028
rect 455506 488016 455512 488028
rect 292908 487988 455512 488016
rect 292908 487976 292914 487988
rect 455506 487976 455512 487988
rect 455564 487976 455570 488028
rect 158254 487908 158260 487960
rect 158312 487948 158318 487960
rect 334066 487948 334072 487960
rect 158312 487920 334072 487948
rect 158312 487908 158318 487920
rect 334066 487908 334072 487920
rect 334124 487908 334130 487960
rect 66898 487840 66904 487892
rect 66956 487880 66962 487892
rect 300118 487880 300124 487892
rect 66956 487852 300124 487880
rect 66956 487840 66962 487852
rect 300118 487840 300124 487852
rect 300176 487840 300182 487892
rect 88242 487772 88248 487824
rect 88300 487812 88306 487824
rect 339494 487812 339500 487824
rect 88300 487784 339500 487812
rect 88300 487772 88306 487784
rect 339494 487772 339500 487784
rect 339552 487772 339558 487824
rect 350534 487772 350540 487824
rect 350592 487812 350598 487824
rect 497458 487812 497464 487824
rect 350592 487784 497464 487812
rect 350592 487772 350598 487784
rect 497458 487772 497464 487784
rect 497516 487772 497522 487824
rect 324498 487160 324504 487212
rect 324556 487200 324562 487212
rect 415118 487200 415124 487212
rect 324556 487172 415124 487200
rect 324556 487160 324562 487172
rect 415118 487160 415124 487172
rect 415176 487200 415182 487212
rect 417878 487200 417884 487212
rect 415176 487172 417884 487200
rect 415176 487160 415182 487172
rect 417878 487160 417884 487172
rect 417936 487160 417942 487212
rect 62758 487092 62764 487144
rect 62816 487132 62822 487144
rect 286318 487132 286324 487144
rect 62816 487104 286324 487132
rect 62816 487092 62822 487104
rect 286318 487092 286324 487104
rect 286376 487092 286382 487144
rect 282914 486616 282920 486668
rect 282972 486656 282978 486668
rect 449894 486656 449900 486668
rect 282972 486628 449900 486656
rect 282972 486616 282978 486628
rect 449894 486616 449900 486628
rect 449952 486616 449958 486668
rect 158162 486548 158168 486600
rect 158220 486588 158226 486600
rect 346486 486588 346492 486600
rect 158220 486560 346492 486588
rect 158220 486548 158226 486560
rect 346486 486548 346492 486560
rect 346544 486548 346550 486600
rect 91002 486480 91008 486532
rect 91060 486520 91066 486532
rect 342346 486520 342352 486532
rect 91060 486492 342352 486520
rect 91060 486480 91066 486492
rect 342346 486480 342352 486492
rect 342404 486480 342410 486532
rect 208578 486412 208584 486464
rect 208636 486452 208642 486464
rect 573358 486452 573364 486464
rect 208636 486424 573364 486452
rect 208636 486412 208642 486424
rect 573358 486412 573364 486424
rect 573416 486412 573422 486464
rect 285674 485868 285680 485920
rect 285732 485908 285738 485920
rect 286318 485908 286324 485920
rect 285732 485880 286324 485908
rect 285732 485868 285738 485880
rect 286318 485868 286324 485880
rect 286376 485868 286382 485920
rect 73982 485732 73988 485784
rect 74040 485772 74046 485784
rect 324498 485772 324504 485784
rect 74040 485744 324504 485772
rect 74040 485732 74046 485744
rect 324498 485732 324504 485744
rect 324556 485732 324562 485784
rect 156782 485188 156788 485240
rect 156840 485228 156846 485240
rect 356054 485228 356060 485240
rect 156840 485200 356060 485228
rect 156840 485188 156846 485200
rect 356054 485188 356060 485200
rect 356112 485188 356118 485240
rect 10318 485120 10324 485172
rect 10376 485160 10382 485172
rect 221090 485160 221096 485172
rect 10376 485132 221096 485160
rect 10376 485120 10382 485132
rect 221090 485120 221096 485132
rect 221148 485120 221154 485172
rect 96522 485052 96528 485104
rect 96580 485092 96586 485104
rect 347774 485092 347780 485104
rect 96580 485064 347780 485092
rect 96580 485052 96586 485064
rect 347774 485052 347780 485064
rect 347832 485052 347838 485104
rect 209038 484372 209044 484424
rect 209096 484412 209102 484424
rect 580166 484412 580172 484424
rect 209096 484384 580172 484412
rect 209096 484372 209102 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 281810 484304 281816 484356
rect 281868 484344 281874 484356
rect 413922 484344 413928 484356
rect 281868 484316 413928 484344
rect 281868 484304 281874 484316
rect 413922 484304 413928 484316
rect 413980 484344 413986 484356
rect 417878 484344 417884 484356
rect 413980 484316 417884 484344
rect 413980 484304 413986 484316
rect 417878 484304 417884 484316
rect 417936 484304 417942 484356
rect 163590 483828 163596 483880
rect 163648 483868 163654 483880
rect 327166 483868 327172 483880
rect 163648 483840 327172 483868
rect 163648 483828 163654 483840
rect 327166 483828 327172 483840
rect 327224 483828 327230 483880
rect 417878 483828 417884 483880
rect 417936 483868 417942 483880
rect 443638 483868 443644 483880
rect 417936 483840 443644 483868
rect 417936 483828 417942 483840
rect 443638 483828 443644 483840
rect 443696 483828 443702 483880
rect 3418 483760 3424 483812
rect 3476 483800 3482 483812
rect 222470 483800 222476 483812
rect 3476 483772 222476 483800
rect 3476 483760 3482 483772
rect 222470 483760 222476 483772
rect 222528 483760 222534 483812
rect 296898 483760 296904 483812
rect 296956 483800 296962 483812
rect 458174 483800 458180 483812
rect 296956 483772 458180 483800
rect 296956 483760 296962 483772
rect 458174 483760 458180 483772
rect 458232 483760 458238 483812
rect 86862 483692 86868 483744
rect 86920 483732 86926 483744
rect 336826 483732 336832 483744
rect 86920 483704 336832 483732
rect 86920 483692 86926 483704
rect 336826 483692 336832 483704
rect 336884 483692 336890 483744
rect 345014 483692 345020 483744
rect 345072 483732 345078 483744
rect 492674 483732 492680 483744
rect 345072 483704 492680 483732
rect 345072 483692 345078 483704
rect 492674 483692 492680 483704
rect 492732 483692 492738 483744
rect 205634 483624 205640 483676
rect 205692 483664 205698 483676
rect 570598 483664 570604 483676
rect 205692 483636 570604 483664
rect 205692 483624 205698 483636
rect 570598 483624 570604 483636
rect 570656 483624 570662 483676
rect 305086 482468 305092 482520
rect 305144 482508 305150 482520
rect 462406 482508 462412 482520
rect 305144 482480 462412 482508
rect 305144 482468 305150 482480
rect 462406 482468 462412 482480
rect 462464 482468 462470 482520
rect 71682 482400 71688 482452
rect 71740 482440 71746 482452
rect 316126 482440 316132 482452
rect 71740 482412 316132 482440
rect 71740 482400 71746 482412
rect 316126 482400 316132 482412
rect 316184 482400 316190 482452
rect 84102 482332 84108 482384
rect 84160 482372 84166 482384
rect 332594 482372 332600 482384
rect 84160 482344 332600 482372
rect 84160 482332 84166 482344
rect 332594 482332 332600 482344
rect 332652 482332 332658 482384
rect 338114 482332 338120 482384
rect 338172 482372 338178 482384
rect 487154 482372 487160 482384
rect 338172 482344 487160 482372
rect 338172 482332 338178 482344
rect 487154 482332 487160 482344
rect 487212 482332 487218 482384
rect 205726 482264 205732 482316
rect 205784 482304 205790 482316
rect 566458 482304 566464 482316
rect 205784 482276 566464 482304
rect 205784 482264 205790 482276
rect 566458 482264 566464 482276
rect 566516 482264 566522 482316
rect 415026 481584 415032 481636
rect 415084 481624 415090 481636
rect 449158 481624 449164 481636
rect 415084 481596 449164 481624
rect 415084 481584 415090 481596
rect 449158 481584 449164 481596
rect 449216 481584 449222 481636
rect 201494 481040 201500 481092
rect 201552 481080 201558 481092
rect 215570 481080 215576 481092
rect 201552 481052 215576 481080
rect 201552 481040 201558 481052
rect 215570 481040 215576 481052
rect 215628 481040 215634 481092
rect 309134 481040 309140 481092
rect 309192 481080 309198 481092
rect 465166 481080 465172 481092
rect 309192 481052 465172 481080
rect 309192 481040 309198 481052
rect 465166 481040 465172 481052
rect 465224 481040 465230 481092
rect 66162 480972 66168 481024
rect 66220 481012 66226 481024
rect 309226 481012 309232 481024
rect 66220 480984 309232 481012
rect 66220 480972 66226 480984
rect 309226 480972 309232 480984
rect 309284 480972 309290 481024
rect 81342 480904 81348 480956
rect 81400 480944 81406 480956
rect 329926 480944 329932 480956
rect 81400 480916 329932 480944
rect 81400 480904 81406 480916
rect 329926 480904 329932 480916
rect 329984 480904 329990 480956
rect 335354 480904 335360 480956
rect 335412 480944 335418 480956
rect 485774 480944 485780 480956
rect 335412 480916 485780 480944
rect 335412 480904 335418 480916
rect 485774 480904 485780 480916
rect 485832 480904 485838 480956
rect 301498 480224 301504 480276
rect 301556 480264 301562 480276
rect 415026 480264 415032 480276
rect 301556 480236 415032 480264
rect 301556 480224 301562 480236
rect 415026 480224 415032 480236
rect 415084 480224 415090 480276
rect 319438 480156 319444 480208
rect 319496 480196 319502 480208
rect 419350 480196 419356 480208
rect 319496 480168 419356 480196
rect 319496 480156 319502 480168
rect 419350 480156 419356 480168
rect 419408 480156 419414 480208
rect 278774 479612 278780 479664
rect 278832 479652 278838 479664
rect 447134 479652 447140 479664
rect 278832 479624 447140 479652
rect 278832 479612 278838 479624
rect 447134 479612 447140 479624
rect 447192 479612 447198 479664
rect 159358 479544 159364 479596
rect 159416 479584 159422 479596
rect 340966 479584 340972 479596
rect 159416 479556 340972 479584
rect 159416 479544 159422 479556
rect 340966 479544 340972 479556
rect 341024 479544 341030 479596
rect 93762 479476 93768 479528
rect 93820 479516 93826 479528
rect 345106 479516 345112 479528
rect 93820 479488 345112 479516
rect 93820 479476 93826 479488
rect 345106 479476 345112 479488
rect 345164 479476 345170 479528
rect 419350 479476 419356 479528
rect 419408 479516 419414 479528
rect 419994 479516 420000 479528
rect 419408 479488 420000 479516
rect 419408 479476 419414 479488
rect 419994 479476 420000 479488
rect 420052 479516 420058 479528
rect 453298 479516 453304 479528
rect 420052 479488 453304 479516
rect 420052 479476 420058 479488
rect 453298 479476 453304 479488
rect 453356 479476 453362 479528
rect 318886 478864 318892 478916
rect 318944 478904 318950 478916
rect 319438 478904 319444 478916
rect 318944 478876 319444 478904
rect 318944 478864 318950 478876
rect 319438 478864 319444 478876
rect 319496 478864 319502 478916
rect 104802 478252 104808 478304
rect 104860 478292 104866 478304
rect 357526 478292 357532 478304
rect 104860 478264 357532 478292
rect 104860 478252 104866 478264
rect 357526 478252 357532 478264
rect 357584 478252 357590 478304
rect 19426 478184 19432 478236
rect 19484 478224 19490 478236
rect 295334 478224 295340 478236
rect 19484 478196 295340 478224
rect 19484 478184 19490 478196
rect 295334 478184 295340 478196
rect 295392 478184 295398 478236
rect 332686 478184 332692 478236
rect 332744 478224 332750 478236
rect 483014 478224 483020 478236
rect 332744 478196 483020 478224
rect 332744 478184 332750 478196
rect 483014 478184 483020 478196
rect 483072 478184 483078 478236
rect 205818 478116 205824 478168
rect 205876 478156 205882 478168
rect 562318 478156 562324 478168
rect 205876 478128 562324 478156
rect 205876 478116 205882 478128
rect 562318 478116 562324 478128
rect 562376 478116 562382 478168
rect 68278 476892 68284 476944
rect 68336 476932 68342 476944
rect 307018 476932 307024 476944
rect 68336 476904 307024 476932
rect 68336 476892 68342 476904
rect 307018 476892 307024 476904
rect 307076 476892 307082 476944
rect 115842 476824 115848 476876
rect 115900 476864 115906 476876
rect 371234 476864 371240 476876
rect 115900 476836 371240 476864
rect 115900 476824 115906 476836
rect 371234 476824 371240 476836
rect 371292 476824 371298 476876
rect 19334 476756 19340 476808
rect 19392 476796 19398 476808
rect 311894 476796 311900 476808
rect 19392 476768 311900 476796
rect 19392 476756 19398 476768
rect 311894 476756 311900 476768
rect 311952 476756 311958 476808
rect 321554 476756 321560 476808
rect 321612 476796 321618 476808
rect 476114 476796 476120 476808
rect 321612 476768 476120 476796
rect 321612 476756 321618 476768
rect 476114 476756 476120 476768
rect 476172 476756 476178 476808
rect 209958 475532 209964 475584
rect 210016 475572 210022 475584
rect 392578 475572 392584 475584
rect 210016 475544 392584 475572
rect 210016 475532 210022 475544
rect 392578 475532 392584 475544
rect 392636 475532 392642 475584
rect 11698 475464 11704 475516
rect 11756 475504 11762 475516
rect 220906 475504 220912 475516
rect 11756 475476 220912 475504
rect 11756 475464 11762 475476
rect 220906 475464 220912 475476
rect 220964 475464 220970 475516
rect 287146 475464 287152 475516
rect 287204 475504 287210 475516
rect 403618 475504 403624 475516
rect 287204 475476 403624 475504
rect 287204 475464 287210 475476
rect 403618 475464 403624 475476
rect 403676 475464 403682 475516
rect 73798 475396 73804 475448
rect 73856 475436 73862 475448
rect 322198 475436 322204 475448
rect 73856 475408 322204 475436
rect 73856 475396 73862 475408
rect 322198 475396 322204 475408
rect 322256 475396 322262 475448
rect 99282 475328 99288 475380
rect 99340 475368 99346 475380
rect 352006 475368 352012 475380
rect 99340 475340 352012 475368
rect 99340 475328 99346 475340
rect 352006 475328 352012 475340
rect 352064 475328 352070 475380
rect 356146 475328 356152 475380
rect 356204 475368 356210 475380
rect 502334 475368 502340 475380
rect 356204 475340 502340 475368
rect 356204 475328 356210 475340
rect 502334 475328 502340 475340
rect 502392 475328 502398 475380
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 80698 474756 80704 474768
rect 3108 474728 80704 474756
rect 3108 474716 3114 474728
rect 80698 474716 80704 474728
rect 80756 474716 80762 474768
rect 303798 474172 303804 474224
rect 303856 474212 303862 474224
rect 417418 474212 417424 474224
rect 303856 474184 417424 474212
rect 303856 474172 303862 474184
rect 417418 474172 417424 474184
rect 417476 474172 417482 474224
rect 43438 474104 43444 474156
rect 43496 474144 43502 474156
rect 290458 474144 290464 474156
rect 43496 474116 290464 474144
rect 43496 474104 43502 474116
rect 290458 474104 290464 474116
rect 290516 474104 290522 474156
rect 294046 474104 294052 474156
rect 294104 474144 294110 474156
rect 414658 474144 414664 474156
rect 294104 474116 414664 474144
rect 294104 474104 294110 474116
rect 414658 474104 414664 474116
rect 414716 474104 414722 474156
rect 114462 474036 114468 474088
rect 114520 474076 114526 474088
rect 368750 474076 368756 474088
rect 114520 474048 368756 474076
rect 114520 474036 114526 474048
rect 368750 474036 368756 474048
rect 368808 474036 368814 474088
rect 379514 474036 379520 474088
rect 379572 474076 379578 474088
rect 523034 474076 523040 474088
rect 379572 474048 523040 474076
rect 379572 474036 379578 474048
rect 523034 474036 523040 474048
rect 523092 474036 523098 474088
rect 205910 473968 205916 474020
rect 205968 474008 205974 474020
rect 558270 474008 558276 474020
rect 205968 473980 558276 474008
rect 205968 473968 205974 473980
rect 558270 473968 558276 473980
rect 558328 473968 558334 474020
rect 405642 473288 405648 473340
rect 405700 473328 405706 473340
rect 406378 473328 406384 473340
rect 405700 473300 406384 473328
rect 405700 473288 405706 473300
rect 406378 473288 406384 473300
rect 406436 473288 406442 473340
rect 162210 472812 162216 472864
rect 162268 472852 162274 472864
rect 324498 472852 324504 472864
rect 162268 472824 324504 472852
rect 162268 472812 162274 472824
rect 324498 472812 324504 472824
rect 324556 472812 324562 472864
rect 158070 472744 158076 472796
rect 158128 472784 158134 472796
rect 353386 472784 353392 472796
rect 158128 472756 353392 472784
rect 158128 472744 158134 472756
rect 353386 472744 353392 472756
rect 353444 472744 353450 472796
rect 76558 472676 76564 472728
rect 76616 472716 76622 472728
rect 331214 472716 331220 472728
rect 76616 472688 331220 472716
rect 76616 472676 76622 472688
rect 331214 472676 331220 472688
rect 331272 472676 331278 472728
rect 17678 472608 17684 472660
rect 17736 472648 17742 472660
rect 308490 472648 308496 472660
rect 17736 472620 308496 472648
rect 17736 472608 17742 472620
rect 308490 472608 308496 472620
rect 308548 472608 308554 472660
rect 358814 472608 358820 472660
rect 358872 472648 358878 472660
rect 504358 472648 504364 472660
rect 358872 472620 504364 472648
rect 358872 472608 358878 472620
rect 504358 472608 504364 472620
rect 504416 472608 504422 472660
rect 311894 471996 311900 472048
rect 311952 472036 311958 472048
rect 405642 472036 405648 472048
rect 311952 472008 405648 472036
rect 311952 471996 311958 472008
rect 405642 471996 405648 472008
rect 405700 471996 405706 472048
rect 75178 471928 75184 471980
rect 75236 471968 75242 471980
rect 328546 471968 328552 471980
rect 75236 471940 328552 471968
rect 75236 471928 75242 471940
rect 328546 471928 328552 471940
rect 328604 471968 328610 471980
rect 329098 471968 329104 471980
rect 328604 471940 329104 471968
rect 328604 471928 328610 471940
rect 329098 471928 329104 471940
rect 329156 471928 329162 471980
rect 414842 471928 414848 471980
rect 414900 471968 414906 471980
rect 457438 471968 457444 471980
rect 414900 471940 457444 471968
rect 414900 471928 414906 471940
rect 457438 471928 457444 471940
rect 457496 471928 457502 471980
rect 166258 471384 166264 471436
rect 166316 471424 166322 471436
rect 219618 471424 219624 471436
rect 166316 471396 219624 471424
rect 166316 471384 166322 471396
rect 219618 471384 219624 471396
rect 219676 471384 219682 471436
rect 331214 471384 331220 471436
rect 331272 471424 331278 471436
rect 414842 471424 414848 471436
rect 331272 471396 414848 471424
rect 331272 471384 331278 471396
rect 414842 471384 414848 471396
rect 414900 471384 414906 471436
rect 166350 471316 166356 471368
rect 166408 471356 166414 471368
rect 343726 471356 343732 471368
rect 166408 471328 343732 471356
rect 166408 471316 166414 471328
rect 343726 471316 343732 471328
rect 343784 471316 343790 471368
rect 53742 471248 53748 471300
rect 53800 471288 53806 471300
rect 288526 471288 288532 471300
rect 53800 471260 288532 471288
rect 53800 471248 53806 471260
rect 288526 471248 288532 471260
rect 288584 471248 288590 471300
rect 311986 471248 311992 471300
rect 312044 471288 312050 471300
rect 467926 471288 467932 471300
rect 312044 471260 467932 471288
rect 312044 471248 312050 471260
rect 467926 471248 467932 471260
rect 467984 471248 467990 471300
rect 204254 470568 204260 470620
rect 204312 470608 204318 470620
rect 579982 470608 579988 470620
rect 204312 470580 579988 470608
rect 204312 470568 204318 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 69658 470500 69664 470552
rect 69716 470540 69722 470552
rect 311158 470540 311164 470552
rect 69716 470512 311164 470540
rect 69716 470500 69722 470512
rect 311158 470500 311164 470512
rect 311216 470500 311222 470552
rect 417694 470500 417700 470552
rect 417752 470540 417758 470552
rect 450538 470540 450544 470552
rect 417752 470512 450544 470540
rect 417752 470500 417758 470512
rect 450538 470500 450544 470512
rect 450596 470500 450602 470552
rect 118602 469888 118608 469940
rect 118660 469928 118666 469940
rect 375374 469928 375380 469940
rect 118660 469900 375380 469928
rect 118660 469888 118666 469900
rect 375374 469888 375380 469900
rect 375432 469888 375438 469940
rect 17586 469820 17592 469872
rect 17644 469860 17650 469872
rect 300762 469860 300768 469872
rect 17644 469832 300768 469860
rect 17644 469820 17650 469832
rect 300762 469820 300768 469832
rect 300820 469820 300826 469872
rect 371326 469820 371332 469872
rect 371384 469860 371390 469872
rect 514754 469860 514760 469872
rect 371384 469832 514760 469860
rect 371384 469820 371390 469832
rect 514754 469820 514760 469832
rect 514812 469820 514818 469872
rect 307018 469344 307024 469396
rect 307076 469384 307082 469396
rect 307076 469356 316034 469384
rect 307076 469344 307082 469356
rect 310514 469276 310520 469328
rect 310572 469316 310578 469328
rect 311158 469316 311164 469328
rect 310572 469288 311164 469316
rect 310572 469276 310578 469288
rect 311158 469276 311164 469288
rect 311216 469276 311222 469328
rect 316006 469316 316034 469356
rect 417694 469316 417700 469328
rect 316006 469288 417700 469316
rect 417694 469276 417700 469288
rect 417752 469276 417758 469328
rect 303706 469208 303712 469260
rect 303764 469248 303770 469260
rect 304350 469248 304356 469260
rect 303764 469220 304356 469248
rect 303764 469208 303770 469220
rect 304350 469208 304356 469220
rect 304408 469248 304414 469260
rect 413922 469248 413928 469260
rect 304408 469220 413928 469248
rect 304408 469208 304414 469220
rect 413922 469208 413928 469220
rect 413980 469248 413986 469260
rect 414566 469248 414572 469260
rect 413980 469220 414572 469248
rect 413980 469208 413986 469220
rect 414566 469208 414572 469220
rect 414624 469208 414630 469260
rect 300762 469140 300768 469192
rect 300820 469180 300826 469192
rect 407850 469180 407856 469192
rect 300820 469152 407856 469180
rect 300820 469140 300826 469152
rect 407850 469140 407856 469152
rect 407908 469140 407914 469192
rect 414750 469140 414756 469192
rect 414808 469180 414814 469192
rect 447778 469180 447784 469192
rect 414808 469152 447784 469180
rect 414808 469140 414814 469152
rect 447778 469140 447784 469152
rect 447836 469140 447842 469192
rect 201310 468664 201316 468716
rect 201368 468704 201374 468716
rect 252646 468704 252652 468716
rect 201368 468676 252652 468704
rect 201368 468664 201374 468676
rect 252646 468664 252652 468676
rect 252704 468664 252710 468716
rect 300118 468664 300124 468716
rect 300176 468704 300182 468716
rect 414566 468704 414572 468716
rect 300176 468676 414572 468704
rect 300176 468664 300182 468676
rect 414566 468664 414572 468676
rect 414624 468704 414630 468716
rect 414750 468704 414756 468716
rect 414624 468676 414756 468704
rect 414624 468664 414630 468676
rect 414750 468664 414756 468676
rect 414808 468664 414814 468716
rect 197262 468596 197268 468648
rect 197320 468636 197326 468648
rect 249978 468636 249984 468648
rect 197320 468608 249984 468636
rect 197320 468596 197326 468608
rect 249978 468596 249984 468608
rect 250036 468596 250042 468648
rect 284478 468596 284484 468648
rect 284536 468636 284542 468648
rect 418798 468636 418804 468648
rect 284536 468608 418804 468636
rect 284536 468596 284542 468608
rect 418798 468596 418804 468608
rect 418856 468596 418862 468648
rect 167638 468528 167644 468580
rect 167696 468568 167702 468580
rect 331306 468568 331312 468580
rect 167696 468540 331312 468568
rect 167696 468528 167702 468540
rect 331306 468528 331312 468540
rect 331364 468528 331370 468580
rect 16850 468460 16856 468512
rect 16908 468500 16914 468512
rect 295426 468500 295432 468512
rect 16908 468472 295432 468500
rect 16908 468460 16914 468472
rect 295426 468460 295432 468472
rect 295484 468460 295490 468512
rect 363046 468460 363052 468512
rect 363104 468500 363110 468512
rect 507854 468500 507860 468512
rect 363104 468472 507860 468500
rect 363104 468460 363110 468472
rect 507854 468460 507860 468472
rect 507912 468460 507918 468512
rect 299474 467848 299480 467900
rect 299532 467888 299538 467900
rect 300118 467888 300124 467900
rect 299532 467860 300124 467888
rect 299532 467848 299538 467860
rect 300118 467848 300124 467860
rect 300176 467848 300182 467900
rect 313366 467236 313372 467288
rect 313424 467276 313430 467288
rect 388438 467276 388444 467288
rect 313424 467248 388444 467276
rect 313424 467236 313430 467248
rect 388438 467236 388444 467248
rect 388496 467236 388502 467288
rect 157978 467168 157984 467220
rect 158036 467208 158042 467220
rect 321646 467208 321652 467220
rect 158036 467180 321652 467208
rect 158036 467168 158042 467180
rect 321646 467168 321652 467180
rect 321704 467168 321710 467220
rect 16666 467100 16672 467152
rect 16724 467140 16730 467152
rect 291286 467140 291292 467152
rect 16724 467112 291292 467140
rect 16724 467100 16730 467112
rect 291286 467100 291292 467112
rect 291344 467100 291350 467152
rect 368566 467100 368572 467152
rect 368624 467140 368630 467152
rect 512638 467140 512644 467152
rect 368624 467112 512644 467140
rect 368624 467100 368630 467112
rect 512638 467100 512644 467112
rect 512696 467100 512702 467152
rect 295426 466488 295432 466540
rect 295484 466528 295490 466540
rect 295484 466500 393314 466528
rect 295484 466488 295490 466500
rect 19058 466420 19064 466472
rect 19116 466460 19122 466472
rect 42794 466460 42800 466472
rect 19116 466432 42800 466460
rect 19116 466420 19122 466432
rect 42794 466420 42800 466432
rect 42852 466460 42858 466472
rect 43622 466460 43628 466472
rect 42852 466432 43628 466460
rect 42852 466420 42858 466432
rect 43622 466420 43628 466432
rect 43680 466420 43686 466472
rect 79410 466420 79416 466472
rect 79468 466460 79474 466472
rect 80054 466460 80060 466472
rect 79468 466432 80060 466460
rect 79468 466420 79474 466432
rect 80054 466420 80060 466432
rect 80112 466460 80118 466472
rect 338298 466460 338304 466472
rect 80112 466432 338304 466460
rect 80112 466420 80118 466432
rect 338298 466420 338304 466432
rect 338356 466460 338362 466472
rect 338758 466460 338764 466472
rect 338356 466432 338764 466460
rect 338356 466420 338362 466432
rect 338758 466420 338764 466432
rect 338816 466420 338822 466472
rect 393286 466460 393314 466500
rect 411162 466460 411168 466472
rect 393286 466432 411168 466460
rect 411162 466420 411168 466432
rect 411220 466460 411226 466472
rect 411898 466460 411904 466472
rect 411220 466432 411904 466460
rect 411220 466420 411226 466432
rect 411898 466420 411904 466432
rect 411956 466420 411962 466472
rect 198642 466352 198648 466404
rect 198700 466392 198706 466404
rect 241698 466392 241704 466404
rect 198700 466364 241704 466392
rect 198700 466352 198706 466364
rect 241698 466352 241704 466364
rect 241756 466352 241762 466404
rect 411254 466352 411260 466404
rect 411312 466392 411318 466404
rect 414934 466392 414940 466404
rect 411312 466364 414940 466392
rect 411312 466352 411318 466364
rect 414934 466352 414940 466364
rect 414992 466392 414998 466404
rect 458818 466392 458824 466404
rect 414992 466364 458824 466392
rect 414992 466352 414998 466364
rect 458818 466352 458824 466364
rect 458876 466352 458882 466404
rect 202414 466284 202420 466336
rect 202472 466324 202478 466336
rect 248506 466324 248512 466336
rect 202472 466296 248512 466324
rect 202472 466284 202478 466296
rect 248506 466284 248512 466296
rect 248564 466284 248570 466336
rect 195698 466216 195704 466268
rect 195756 466256 195762 466268
rect 243078 466256 243084 466268
rect 195756 466228 243084 466256
rect 195756 466216 195762 466228
rect 243078 466216 243084 466228
rect 243136 466216 243142 466268
rect 199378 466148 199384 466200
rect 199436 466188 199442 466200
rect 247218 466188 247224 466200
rect 199436 466160 247224 466188
rect 199436 466148 199442 466160
rect 247218 466148 247224 466160
rect 247276 466148 247282 466200
rect 195606 466080 195612 466132
rect 195664 466120 195670 466132
rect 245838 466120 245844 466132
rect 195664 466092 245844 466120
rect 195664 466080 195670 466092
rect 245838 466080 245844 466092
rect 245896 466080 245902 466132
rect 202322 466012 202328 466064
rect 202380 466052 202386 466064
rect 252738 466052 252744 466064
rect 202380 466024 252744 466052
rect 202380 466012 202386 466024
rect 252738 466012 252744 466024
rect 252796 466012 252802 466064
rect 198550 465944 198556 465996
rect 198608 465984 198614 465996
rect 251358 465984 251364 465996
rect 198608 465956 251364 465984
rect 198608 465944 198614 465956
rect 251358 465944 251364 465956
rect 251416 465944 251422 465996
rect 195790 465876 195796 465928
rect 195848 465916 195854 465928
rect 250070 465916 250076 465928
rect 195848 465888 250076 465916
rect 195848 465876 195854 465888
rect 250070 465876 250076 465888
rect 250128 465876 250134 465928
rect 197906 465808 197912 465860
rect 197964 465848 197970 465860
rect 310606 465848 310612 465860
rect 197964 465820 310612 465848
rect 197964 465808 197970 465820
rect 310606 465808 310612 465820
rect 310664 465808 310670 465860
rect 43622 465740 43628 465792
rect 43680 465780 43686 465792
rect 281718 465780 281724 465792
rect 43680 465752 281724 465780
rect 43680 465740 43686 465752
rect 281718 465740 281724 465752
rect 281776 465740 281782 465792
rect 301498 465740 301504 465792
rect 301556 465780 301562 465792
rect 304258 465780 304264 465792
rect 301556 465752 304264 465780
rect 301556 465740 301562 465752
rect 304258 465740 304264 465752
rect 304316 465740 304322 465792
rect 365898 465740 365904 465792
rect 365956 465780 365962 465792
rect 510614 465780 510620 465792
rect 365956 465752 510620 465780
rect 365956 465740 365962 465752
rect 510614 465740 510620 465752
rect 510672 465740 510678 465792
rect 126882 465672 126888 465724
rect 126940 465712 126946 465724
rect 383654 465712 383660 465724
rect 126940 465684 383660 465712
rect 126940 465672 126946 465684
rect 383654 465672 383660 465684
rect 383712 465672 383718 465724
rect 201402 465604 201408 465656
rect 201460 465644 201466 465656
rect 240318 465644 240324 465656
rect 201460 465616 240324 465644
rect 201460 465604 201466 465616
rect 240318 465604 240324 465616
rect 240376 465604 240382 465656
rect 65518 465536 65524 465588
rect 65576 465576 65582 465588
rect 66254 465576 66260 465588
rect 65576 465548 66260 465576
rect 65576 465536 65582 465548
rect 66254 465536 66260 465548
rect 66312 465536 66318 465588
rect 199286 465536 199292 465588
rect 199344 465576 199350 465588
rect 237466 465576 237472 465588
rect 199344 465548 237472 465576
rect 199344 465536 199350 465548
rect 237466 465536 237472 465548
rect 237524 465536 237530 465588
rect 409782 465536 409788 465588
rect 409840 465576 409846 465588
rect 410610 465576 410616 465588
rect 409840 465548 410616 465576
rect 409840 465536 409846 465548
rect 410610 465536 410616 465548
rect 410668 465536 410674 465588
rect 291286 465128 291292 465180
rect 291344 465168 291350 465180
rect 409782 465168 409788 465180
rect 291344 465140 409788 465168
rect 291344 465128 291350 465140
rect 409782 465128 409788 465140
rect 409840 465128 409846 465180
rect 18966 465060 18972 465112
rect 19024 465100 19030 465112
rect 38654 465100 38660 465112
rect 19024 465072 38660 465100
rect 19024 465060 19030 465072
rect 38654 465060 38660 465072
rect 38712 465100 38718 465112
rect 38712 465072 39988 465100
rect 38712 465060 38718 465072
rect 39960 465032 39988 465072
rect 66254 465060 66260 465112
rect 66312 465100 66318 465112
rect 295702 465100 295708 465112
rect 66312 465072 295708 465100
rect 66312 465060 66318 465072
rect 295702 465060 295708 465072
rect 295760 465060 295766 465112
rect 336642 465060 336648 465112
rect 336700 465100 336706 465112
rect 411254 465100 411260 465112
rect 336700 465072 411260 465100
rect 336700 465060 336706 465072
rect 411254 465060 411260 465072
rect 411312 465100 411318 465112
rect 412542 465100 412548 465112
rect 411312 465072 412548 465100
rect 411312 465060 411318 465072
rect 412542 465060 412548 465072
rect 412600 465060 412606 465112
rect 277486 465032 277492 465044
rect 39960 465004 277492 465032
rect 277486 464992 277492 465004
rect 277544 465032 277550 465044
rect 278038 465032 278044 465044
rect 277544 465004 278044 465032
rect 277544 464992 277550 465004
rect 278038 464992 278044 465004
rect 278096 464992 278102 465044
rect 287698 464992 287704 465044
rect 287756 465032 287762 465044
rect 288342 465032 288348 465044
rect 287756 465004 288348 465032
rect 287756 464992 287762 465004
rect 288342 464992 288348 465004
rect 288400 465032 288406 465044
rect 415854 465032 415860 465044
rect 288400 465004 415860 465032
rect 288400 464992 288406 465004
rect 415854 464992 415860 465004
rect 415912 464992 415918 465044
rect 417418 464992 417424 465044
rect 417476 465032 417482 465044
rect 440234 465032 440240 465044
rect 417476 465004 440240 465032
rect 417476 464992 417482 465004
rect 440234 464992 440240 465004
rect 440292 464992 440298 465044
rect 79318 464924 79324 464976
rect 79376 464964 79382 464976
rect 80146 464964 80152 464976
rect 79376 464936 80152 464964
rect 79376 464924 79382 464936
rect 80146 464924 80152 464936
rect 80204 464924 80210 464976
rect 187602 464448 187608 464500
rect 187660 464488 187666 464500
rect 232682 464488 232688 464500
rect 187660 464460 232688 464488
rect 187660 464448 187666 464460
rect 232682 464448 232688 464460
rect 232740 464448 232746 464500
rect 290458 464448 290464 464500
rect 290516 464488 290522 464500
rect 417418 464488 417424 464500
rect 290516 464460 417424 464488
rect 290516 464448 290522 464460
rect 417418 464448 417424 464460
rect 417476 464448 417482 464500
rect 186866 464380 186872 464432
rect 186924 464420 186930 464432
rect 232774 464420 232780 464432
rect 186924 464392 232780 464420
rect 186924 464380 186930 464392
rect 232774 464380 232780 464392
rect 232832 464380 232838 464432
rect 373994 464380 374000 464432
rect 374052 464420 374058 464432
rect 517514 464420 517520 464432
rect 374052 464392 517520 464420
rect 374052 464380 374058 464392
rect 517514 464380 517520 464392
rect 517572 464380 517578 464432
rect 124122 464312 124128 464364
rect 124180 464352 124186 464364
rect 380986 464352 380992 464364
rect 124180 464324 380992 464352
rect 124180 464312 124186 464324
rect 380986 464312 380992 464324
rect 381044 464312 381050 464364
rect 188982 464244 188988 464296
rect 189040 464284 189046 464296
rect 235350 464284 235356 464296
rect 189040 464256 235356 464284
rect 189040 464244 189046 464256
rect 235350 464244 235356 464256
rect 235408 464244 235414 464296
rect 191466 464176 191472 464228
rect 191524 464216 191530 464228
rect 273346 464216 273352 464228
rect 191524 464188 273352 464216
rect 191524 464176 191530 464188
rect 273346 464176 273352 464188
rect 273404 464176 273410 464228
rect 289814 464176 289820 464228
rect 289872 464216 289878 464228
rect 290458 464216 290464 464228
rect 289872 464188 290464 464216
rect 289872 464176 289878 464188
rect 290458 464176 290464 464188
rect 290516 464176 290522 464228
rect 188154 464108 188160 464160
rect 188212 464148 188218 464160
rect 271874 464148 271880 464160
rect 188212 464120 271880 464148
rect 188212 464108 188218 464120
rect 271874 464108 271880 464120
rect 271932 464108 271938 464160
rect 186774 464040 186780 464092
rect 186832 464080 186838 464092
rect 271966 464080 271972 464092
rect 186832 464052 271972 464080
rect 186832 464040 186838 464052
rect 271966 464040 271972 464052
rect 272024 464040 272030 464092
rect 183462 463972 183468 464024
rect 183520 464012 183526 464024
rect 270770 464012 270776 464024
rect 183520 463984 270776 464012
rect 183520 463972 183526 463984
rect 270770 463972 270776 463984
rect 270828 463972 270834 464024
rect 186222 463904 186228 463956
rect 186280 463944 186286 463956
rect 274726 463944 274732 463956
rect 186280 463916 274732 463944
rect 186280 463904 186286 463916
rect 274726 463904 274732 463916
rect 274784 463904 274790 463956
rect 184842 463836 184848 463888
rect 184900 463876 184906 463888
rect 274818 463876 274824 463888
rect 184900 463848 274824 463876
rect 184900 463836 184906 463848
rect 274818 463836 274824 463848
rect 274876 463836 274882 463888
rect 186130 463768 186136 463820
rect 186188 463808 186194 463820
rect 276198 463808 276204 463820
rect 186188 463780 276204 463808
rect 186188 463768 186194 463780
rect 276198 463768 276204 463780
rect 276256 463768 276262 463820
rect 18874 463700 18880 463752
rect 18932 463740 18938 463752
rect 44174 463740 44180 463752
rect 18932 463712 44180 463740
rect 18932 463700 18938 463712
rect 44174 463700 44180 463712
rect 44232 463740 44238 463752
rect 44634 463740 44640 463752
rect 44232 463712 44640 463740
rect 44232 463700 44238 463712
rect 44634 463700 44640 463712
rect 44692 463700 44698 463752
rect 80146 463700 80152 463752
rect 80204 463740 80210 463752
rect 335446 463740 335452 463752
rect 80204 463712 335452 463740
rect 80204 463700 80210 463712
rect 335446 463700 335452 463712
rect 335504 463740 335510 463752
rect 336642 463740 336648 463752
rect 335504 463712 336648 463740
rect 335504 463700 335510 463712
rect 336642 463700 336648 463712
rect 336700 463700 336706 463752
rect 199746 463632 199752 463684
rect 199804 463672 199810 463684
rect 241790 463672 241796 463684
rect 199804 463644 241796 463672
rect 199804 463632 199810 463644
rect 241790 463632 241796 463644
rect 241848 463632 241854 463684
rect 308490 463632 308496 463684
rect 308548 463672 308554 463684
rect 309042 463672 309048 463684
rect 308548 463644 309048 463672
rect 308548 463632 308554 463644
rect 309042 463632 309048 463644
rect 309100 463672 309106 463684
rect 383010 463672 383016 463684
rect 309100 463644 383016 463672
rect 309100 463632 309106 463644
rect 383010 463632 383016 463644
rect 383068 463632 383074 463684
rect 199930 463564 199936 463616
rect 199988 463604 199994 463616
rect 243170 463604 243176 463616
rect 199988 463576 243176 463604
rect 199988 463564 199994 463576
rect 243170 463564 243176 463576
rect 243228 463564 243234 463616
rect 199654 463496 199660 463548
rect 199712 463536 199718 463548
rect 244550 463536 244556 463548
rect 199712 463508 244556 463536
rect 199712 463496 199718 463508
rect 244550 463496 244556 463508
rect 244608 463496 244614 463548
rect 199838 463428 199844 463480
rect 199896 463468 199902 463480
rect 247310 463468 247316 463480
rect 199896 463440 247316 463468
rect 199896 463428 199902 463440
rect 247310 463428 247316 463440
rect 247368 463428 247374 463480
rect 195882 463360 195888 463412
rect 195940 463400 195946 463412
rect 254118 463400 254124 463412
rect 195940 463372 254124 463400
rect 195940 463360 195946 463372
rect 254118 463360 254124 463372
rect 254176 463360 254182 463412
rect 200574 463292 200580 463344
rect 200632 463332 200638 463344
rect 281626 463332 281632 463344
rect 200632 463304 281632 463332
rect 200632 463292 200638 463304
rect 281626 463292 281632 463304
rect 281684 463292 281690 463344
rect 200666 463224 200672 463276
rect 200724 463264 200730 463276
rect 285766 463264 285772 463276
rect 200724 463236 285772 463264
rect 200724 463224 200730 463236
rect 285766 463224 285772 463236
rect 285824 463224 285830 463276
rect 200942 463156 200948 463208
rect 201000 463196 201006 463208
rect 361574 463196 361580 463208
rect 201000 463168 361580 463196
rect 201000 463156 201006 463168
rect 361574 463156 361580 463168
rect 361632 463156 361638 463208
rect 201034 463088 201040 463140
rect 201092 463128 201098 463140
rect 364334 463128 364340 463140
rect 201092 463100 364340 463128
rect 201092 463088 201098 463100
rect 364334 463088 364340 463100
rect 364392 463088 364398 463140
rect 419442 463088 419448 463140
rect 419500 463128 419506 463140
rect 436186 463128 436192 463140
rect 419500 463100 436192 463128
rect 419500 463088 419506 463100
rect 436186 463088 436192 463100
rect 436244 463088 436250 463140
rect 44634 463020 44640 463072
rect 44692 463060 44698 463072
rect 285858 463060 285864 463072
rect 44692 463032 285864 463060
rect 44692 463020 44698 463032
rect 285858 463020 285864 463032
rect 285916 463020 285922 463072
rect 376754 463020 376760 463072
rect 376812 463060 376818 463072
rect 519538 463060 519544 463072
rect 376812 463032 519544 463060
rect 376812 463020 376818 463032
rect 519538 463020 519544 463032
rect 519596 463020 519602 463072
rect 121362 462952 121368 463004
rect 121420 462992 121426 463004
rect 378226 462992 378232 463004
rect 121420 462964 378232 462992
rect 121420 462952 121426 462964
rect 378226 462952 378232 462964
rect 378284 462952 378290 463004
rect 414750 462952 414756 463004
rect 414808 462992 414814 463004
rect 445754 462992 445760 463004
rect 414808 462964 445760 462992
rect 414808 462952 414814 462964
rect 445754 462952 445760 462964
rect 445812 462952 445818 463004
rect 199562 462884 199568 462936
rect 199620 462924 199626 462936
rect 239030 462924 239036 462936
rect 199620 462896 239036 462924
rect 199620 462884 199626 462896
rect 239030 462884 239036 462896
rect 239088 462884 239094 462936
rect 199470 462816 199476 462868
rect 199528 462856 199534 462868
rect 236178 462856 236184 462868
rect 199528 462828 236184 462856
rect 199528 462816 199534 462828
rect 236178 462816 236184 462828
rect 236236 462816 236242 462868
rect 295702 462408 295708 462460
rect 295760 462448 295766 462460
rect 414750 462448 414756 462460
rect 295760 462420 414756 462448
rect 295760 462408 295766 462420
rect 414750 462408 414756 462420
rect 414808 462408 414814 462460
rect 3418 462340 3424 462392
rect 3476 462380 3482 462392
rect 218054 462380 218060 462392
rect 3476 462352 218060 462380
rect 3476 462340 3482 462352
rect 218054 462340 218060 462352
rect 218112 462340 218118 462392
rect 281718 462340 281724 462392
rect 281776 462380 281782 462392
rect 419442 462380 419448 462392
rect 281776 462352 419448 462380
rect 281776 462340 281782 462352
rect 419442 462340 419448 462352
rect 419500 462340 419506 462392
rect 192478 461932 192484 461984
rect 192536 461972 192542 461984
rect 218146 461972 218152 461984
rect 192536 461944 218152 461972
rect 192536 461932 192542 461944
rect 218146 461932 218152 461944
rect 218204 461932 218210 461984
rect 191098 461864 191104 461916
rect 191156 461904 191162 461916
rect 216766 461904 216772 461916
rect 191156 461876 216772 461904
rect 191156 461864 191162 461876
rect 216766 461864 216772 461876
rect 216824 461864 216830 461916
rect 169754 461796 169760 461848
rect 169812 461836 169818 461848
rect 216858 461836 216864 461848
rect 169812 461808 216864 461836
rect 169812 461796 169818 461808
rect 216858 461796 216864 461808
rect 216916 461796 216922 461848
rect 218054 461796 218060 461848
rect 218112 461836 218118 461848
rect 225046 461836 225052 461848
rect 218112 461808 225052 461836
rect 218112 461796 218118 461808
rect 225046 461796 225052 461808
rect 225104 461796 225110 461848
rect 200850 461728 200856 461780
rect 200908 461768 200914 461780
rect 374086 461768 374092 461780
rect 200908 461740 374092 461768
rect 200908 461728 200914 461740
rect 374086 461728 374092 461740
rect 374144 461728 374150 461780
rect 14458 461660 14464 461712
rect 14516 461700 14522 461712
rect 219710 461700 219716 461712
rect 14516 461672 219716 461700
rect 14516 461660 14522 461672
rect 219710 461660 219716 461672
rect 219768 461660 219774 461712
rect 298278 461660 298284 461712
rect 298336 461700 298342 461712
rect 380158 461700 380164 461712
rect 298336 461672 380164 461700
rect 298336 461660 298342 461672
rect 380158 461660 380164 461672
rect 380216 461660 380222 461712
rect 10410 461592 10416 461644
rect 10468 461632 10474 461644
rect 222286 461632 222292 461644
rect 10468 461604 222292 461632
rect 10468 461592 10474 461604
rect 222286 461592 222292 461604
rect 222344 461592 222350 461644
rect 347866 461592 347872 461644
rect 347924 461632 347930 461644
rect 494698 461632 494704 461644
rect 347924 461604 494704 461632
rect 347924 461592 347930 461604
rect 494698 461592 494704 461604
rect 494756 461592 494762 461644
rect 191742 461388 191748 461440
rect 191800 461428 191806 461440
rect 270586 461428 270592 461440
rect 191800 461400 270592 461428
rect 191800 461388 191806 461400
rect 270586 461388 270592 461400
rect 270644 461388 270650 461440
rect 185854 461320 185860 461372
rect 185912 461360 185918 461372
rect 266354 461360 266360 461372
rect 185912 461332 266360 461360
rect 185912 461320 185918 461332
rect 266354 461320 266360 461332
rect 266412 461320 266418 461372
rect 189534 461252 189540 461304
rect 189592 461292 189598 461304
rect 270678 461292 270684 461304
rect 189592 461264 270684 461292
rect 189592 461252 189598 461264
rect 270678 461252 270684 461264
rect 270736 461252 270742 461304
rect 190362 461184 190368 461236
rect 190420 461224 190426 461236
rect 272058 461224 272064 461236
rect 190420 461196 272064 461224
rect 190420 461184 190426 461196
rect 272058 461184 272064 461196
rect 272116 461184 272122 461236
rect 185762 461116 185768 461168
rect 185820 461156 185826 461168
rect 267734 461156 267740 461168
rect 185820 461128 267740 461156
rect 185820 461116 185826 461128
rect 267734 461116 267740 461128
rect 267792 461116 267798 461168
rect 173618 461048 173624 461100
rect 173676 461088 173682 461100
rect 294138 461088 294144 461100
rect 173676 461060 294144 461088
rect 173676 461048 173682 461060
rect 294138 461048 294144 461060
rect 294196 461048 294202 461100
rect 173434 460980 173440 461032
rect 173492 461020 173498 461032
rect 306374 461020 306380 461032
rect 173492 460992 306380 461020
rect 173492 460980 173498 460992
rect 306374 460980 306380 460992
rect 306432 460980 306438 461032
rect 198734 460912 198740 460964
rect 198792 460952 198798 460964
rect 580626 460952 580632 460964
rect 198792 460924 580632 460952
rect 198792 460912 198798 460924
rect 580626 460912 580632 460924
rect 580684 460912 580690 460964
rect 385770 460844 385776 460896
rect 385828 460884 385834 460896
rect 387058 460884 387064 460896
rect 385828 460856 387064 460884
rect 385828 460844 385834 460856
rect 387058 460844 387064 460856
rect 387116 460844 387122 460896
rect 200022 460640 200028 460692
rect 200080 460680 200086 460692
rect 237926 460680 237932 460692
rect 200080 460652 237932 460680
rect 200080 460640 200086 460652
rect 237926 460640 237932 460652
rect 237984 460640 237990 460692
rect 198090 460572 198096 460624
rect 198148 460612 198154 460624
rect 290182 460612 290188 460624
rect 198148 460584 290188 460612
rect 198148 460572 198154 460584
rect 290182 460572 290188 460584
rect 290240 460572 290246 460624
rect 197998 460504 198004 460556
rect 198056 460544 198062 460556
rect 294598 460544 294604 460556
rect 198056 460516 294604 460544
rect 198056 460504 198062 460516
rect 294598 460504 294604 460516
rect 294656 460504 294662 460556
rect 198366 460436 198372 460488
rect 198424 460476 198430 460488
rect 299014 460476 299020 460488
rect 198424 460448 299020 460476
rect 198424 460436 198430 460448
rect 299014 460436 299020 460448
rect 299072 460436 299078 460488
rect 198274 460368 198280 460420
rect 198332 460408 198338 460420
rect 303062 460408 303068 460420
rect 198332 460380 303068 460408
rect 198332 460368 198338 460380
rect 303062 460368 303068 460380
rect 303120 460368 303126 460420
rect 198182 460300 198188 460352
rect 198240 460340 198246 460352
rect 307110 460340 307116 460352
rect 198240 460312 307116 460340
rect 198240 460300 198246 460312
rect 307110 460300 307116 460312
rect 307168 460300 307174 460352
rect 156598 460232 156604 460284
rect 156656 460272 156662 460284
rect 358906 460272 358912 460284
rect 156656 460244 358912 460272
rect 156656 460232 156662 460244
rect 358906 460232 358912 460244
rect 358964 460232 358970 460284
rect 3602 460164 3608 460216
rect 3660 460204 3666 460216
rect 223942 460204 223948 460216
rect 3660 460176 223948 460204
rect 3660 460164 3666 460176
rect 223942 460164 223948 460176
rect 224000 460164 224006 460216
rect 185946 459892 185952 459944
rect 186004 459932 186010 459944
rect 269114 459932 269120 459944
rect 186004 459904 269120 459932
rect 186004 459892 186010 459904
rect 269114 459892 269120 459904
rect 269172 459892 269178 459944
rect 186038 459824 186044 459876
rect 186096 459864 186102 459876
rect 276106 459864 276112 459876
rect 186096 459836 276112 459864
rect 186096 459824 186102 459836
rect 276106 459824 276112 459836
rect 276164 459824 276170 459876
rect 181438 459756 181444 459808
rect 181496 459796 181502 459808
rect 280982 459796 280988 459808
rect 181496 459768 280988 459796
rect 181496 459756 181502 459768
rect 280982 459756 280988 459768
rect 281040 459756 281046 459808
rect 181714 459688 181720 459740
rect 181772 459728 181778 459740
rect 301222 459728 301228 459740
rect 181772 459700 301228 459728
rect 181772 459688 181778 459700
rect 301222 459688 301228 459700
rect 301280 459688 301286 459740
rect 179046 459620 179052 459672
rect 179104 459660 179110 459672
rect 324314 459660 324320 459672
rect 179104 459632 324320 459660
rect 179104 459620 179110 459632
rect 324314 459620 324320 459632
rect 324372 459620 324378 459672
rect 181622 459552 181628 459604
rect 181680 459592 181686 459604
rect 381078 459592 381084 459604
rect 181680 459564 381084 459592
rect 181680 459552 181686 459564
rect 381078 459552 381084 459564
rect 381136 459552 381142 459604
rect 373994 459484 374000 459536
rect 374052 459524 374058 459536
rect 374454 459524 374460 459536
rect 374052 459496 374460 459524
rect 374052 459484 374058 459496
rect 374454 459484 374460 459496
rect 374512 459484 374518 459536
rect 181530 459212 181536 459264
rect 181588 459252 181594 459264
rect 321094 459252 321100 459264
rect 181588 459224 321100 459252
rect 181588 459212 181594 459224
rect 321094 459212 321100 459224
rect 321152 459212 321158 459264
rect 178770 459144 178776 459196
rect 178828 459184 178834 459196
rect 327718 459184 327724 459196
rect 178828 459156 327724 459184
rect 178828 459144 178834 459156
rect 327718 459144 327724 459156
rect 327776 459144 327782 459196
rect 180058 459076 180064 459128
rect 180116 459116 180122 459128
rect 218422 459116 218428 459128
rect 180116 459088 218428 459116
rect 180116 459076 180122 459088
rect 218422 459076 218428 459088
rect 218480 459076 218486 459128
rect 163498 459008 163504 459060
rect 163556 459048 163562 459060
rect 216674 459048 216680 459060
rect 163556 459020 216680 459048
rect 163556 459008 163562 459020
rect 216674 459008 216680 459020
rect 216732 459008 216738 459060
rect 188614 458940 188620 458992
rect 188672 458980 188678 458992
rect 262950 458980 262956 458992
rect 188672 458952 262956 458980
rect 188672 458940 188678 458952
rect 262950 458940 262956 458952
rect 263008 458940 263014 458992
rect 15746 458872 15752 458924
rect 15804 458912 15810 458924
rect 223666 458912 223672 458924
rect 15804 458884 223672 458912
rect 15804 458872 15810 458884
rect 223666 458872 223672 458884
rect 223724 458872 223730 458924
rect 7650 458804 7656 458856
rect 7708 458844 7714 458856
rect 222470 458844 222476 458856
rect 7708 458816 222476 458844
rect 7708 458804 7714 458816
rect 222470 458804 222476 458816
rect 222528 458804 222534 458856
rect 190270 458736 190276 458788
rect 190328 458776 190334 458788
rect 266998 458776 267004 458788
rect 190328 458748 267004 458776
rect 190328 458736 190334 458748
rect 266998 458736 267004 458748
rect 267056 458736 267062 458788
rect 306006 458736 306012 458788
rect 306064 458776 306070 458788
rect 402238 458776 402244 458788
rect 306064 458748 402244 458776
rect 306064 458736 306070 458748
rect 402238 458736 402244 458748
rect 402296 458736 402302 458788
rect 184750 458668 184756 458720
rect 184808 458708 184814 458720
rect 277578 458708 277584 458720
rect 184808 458680 277584 458708
rect 184808 458668 184814 458680
rect 277578 458668 277584 458680
rect 277636 458668 277642 458720
rect 302510 458668 302516 458720
rect 302568 458708 302574 458720
rect 402330 458708 402336 458720
rect 302568 458680 402336 458708
rect 302568 458668 302574 458680
rect 402330 458668 402336 458680
rect 402388 458668 402394 458720
rect 310054 458600 310060 458652
rect 310112 458640 310118 458652
rect 399662 458640 399668 458652
rect 310112 458612 399668 458640
rect 310112 458600 310118 458612
rect 399662 458600 399668 458612
rect 399720 458600 399726 458652
rect 313734 458532 313740 458584
rect 313792 458572 313798 458584
rect 399478 458572 399484 458584
rect 313792 458544 399484 458572
rect 313792 458532 313798 458544
rect 399478 458532 399484 458544
rect 399536 458532 399542 458584
rect 181898 458464 181904 458516
rect 181956 458504 181962 458516
rect 313182 458504 313188 458516
rect 181956 458476 313188 458504
rect 181956 458464 181962 458476
rect 313182 458464 313188 458476
rect 313240 458464 313246 458516
rect 317046 458464 317052 458516
rect 317104 458504 317110 458516
rect 399570 458504 399576 458516
rect 317104 458476 399576 458504
rect 317104 458464 317110 458476
rect 399570 458464 399576 458476
rect 399628 458464 399634 458516
rect 178678 458396 178684 458448
rect 178736 458436 178742 458448
rect 334342 458436 334348 458448
rect 178736 458408 334348 458436
rect 178736 458396 178742 458408
rect 334342 458396 334348 458408
rect 334400 458396 334406 458448
rect 178862 458328 178868 458380
rect 178920 458368 178926 458380
rect 341058 458368 341064 458380
rect 178920 458340 341064 458368
rect 178920 458328 178926 458340
rect 341058 458328 341064 458340
rect 341116 458328 341122 458380
rect 198826 458260 198832 458312
rect 198884 458300 198890 458312
rect 580442 458300 580448 458312
rect 198884 458272 580448 458300
rect 198884 458260 198890 458272
rect 580442 458260 580448 458272
rect 580500 458260 580506 458312
rect 199286 458192 199292 458244
rect 199344 458232 199350 458244
rect 580718 458232 580724 458244
rect 199344 458204 580724 458232
rect 199344 458192 199350 458204
rect 580718 458192 580724 458204
rect 580776 458192 580782 458244
rect 80698 457784 80704 457836
rect 80756 457824 80762 457836
rect 224310 457824 224316 457836
rect 80756 457796 224316 457824
rect 80756 457784 80762 457796
rect 224310 457784 224316 457796
rect 224368 457784 224374 457836
rect 353294 457784 353300 457836
rect 353352 457824 353358 457836
rect 353846 457824 353852 457836
rect 353352 457796 353852 457824
rect 353352 457784 353358 457796
rect 353846 457784 353852 457796
rect 353904 457784 353910 457836
rect 210050 457716 210056 457768
rect 210108 457756 210114 457768
rect 400858 457756 400864 457768
rect 210108 457728 400864 457756
rect 210108 457716 210114 457728
rect 400858 457716 400864 457728
rect 400916 457716 400922 457768
rect 14550 457648 14556 457700
rect 14608 457688 14614 457700
rect 220998 457688 221004 457700
rect 14608 457660 221004 457688
rect 14608 457648 14614 457660
rect 220998 457648 221004 457660
rect 221056 457648 221062 457700
rect 4798 457580 4804 457632
rect 4856 457620 4862 457632
rect 220814 457620 220820 457632
rect 4856 457592 220820 457620
rect 4856 457580 4862 457592
rect 220814 457580 220820 457592
rect 220872 457580 220878 457632
rect 208854 457512 208860 457564
rect 208912 457552 208918 457564
rect 565078 457552 565084 457564
rect 208912 457524 565084 457552
rect 208912 457512 208918 457524
rect 565078 457512 565084 457524
rect 565136 457512 565142 457564
rect 207750 457444 207756 457496
rect 207808 457484 207814 457496
rect 563698 457484 563704 457496
rect 207808 457456 563704 457484
rect 207808 457444 207814 457456
rect 563698 457444 563704 457456
rect 563756 457444 563762 457496
rect 201494 457308 201500 457360
rect 201552 457348 201558 457360
rect 209130 457348 209136 457360
rect 201552 457320 209136 457348
rect 201552 457308 201558 457320
rect 209130 457308 209136 457320
rect 209188 457308 209194 457360
rect 191650 457240 191656 457292
rect 191708 457280 191714 457292
rect 264974 457280 264980 457292
rect 191708 457252 264980 457280
rect 191708 457240 191714 457252
rect 264974 457240 264980 457252
rect 265032 457240 265038 457292
rect 186958 457172 186964 457224
rect 187016 457212 187022 457224
rect 319622 457212 319628 457224
rect 187016 457184 319628 457212
rect 187016 457172 187022 457184
rect 319622 457172 319628 457184
rect 319680 457172 319686 457224
rect 187050 457104 187056 457156
rect 187108 457144 187114 457156
rect 326246 457144 326252 457156
rect 187108 457116 326252 457144
rect 187108 457104 187114 457116
rect 326246 457104 326252 457116
rect 326304 457104 326310 457156
rect 184198 457036 184204 457088
rect 184256 457076 184262 457088
rect 360194 457076 360200 457088
rect 184256 457048 360200 457076
rect 184256 457036 184262 457048
rect 360194 457036 360200 457048
rect 360252 457036 360258 457088
rect 184290 456968 184296 457020
rect 184348 457008 184354 457020
rect 365990 457008 365996 457020
rect 184348 456980 365996 457008
rect 184348 456968 184354 456980
rect 365990 456968 365996 456980
rect 366048 456968 366054 457020
rect 204346 456900 204352 456952
rect 204404 456940 204410 456952
rect 394142 456940 394148 456952
rect 204404 456912 394148 456940
rect 204404 456900 204410 456912
rect 394142 456900 394148 456912
rect 394200 456900 394206 456952
rect 203058 456832 203064 456884
rect 203116 456872 203122 456884
rect 399754 456872 399760 456884
rect 203116 456844 399760 456872
rect 203116 456832 203122 456844
rect 399754 456832 399760 456844
rect 399812 456832 399818 456884
rect 204806 456764 204812 456816
rect 204864 456804 204870 456816
rect 209038 456804 209044 456816
rect 204864 456776 209044 456804
rect 204864 456764 204870 456776
rect 209038 456764 209044 456776
rect 209096 456764 209102 456816
rect 209130 456764 209136 456816
rect 209188 456804 209194 456816
rect 403618 456804 403624 456816
rect 209188 456776 403624 456804
rect 209188 456764 209194 456776
rect 403618 456764 403624 456776
rect 403676 456764 403682 456816
rect 200666 456424 200672 456476
rect 200724 456464 200730 456476
rect 209498 456464 209504 456476
rect 200724 456436 209504 456464
rect 200724 456424 200730 456436
rect 209498 456424 209504 456436
rect 209556 456424 209562 456476
rect 181990 456356 181996 456408
rect 182048 456396 182054 456408
rect 293034 456396 293040 456408
rect 182048 456368 293040 456396
rect 182048 456356 182054 456368
rect 293034 456356 293040 456368
rect 293092 456356 293098 456408
rect 183370 456288 183376 456340
rect 183428 456328 183434 456340
rect 269942 456328 269948 456340
rect 183428 456300 269948 456328
rect 183428 456288 183434 456300
rect 269942 456288 269948 456300
rect 270000 456288 270006 456340
rect 310514 456288 310520 456340
rect 310572 456328 310578 456340
rect 311526 456328 311532 456340
rect 310572 456300 311532 456328
rect 310572 456288 310578 456300
rect 311526 456288 311532 456300
rect 311584 456288 311590 456340
rect 322198 456288 322204 456340
rect 322256 456328 322262 456340
rect 419626 456328 419632 456340
rect 322256 456300 419632 456328
rect 322256 456288 322262 456300
rect 419626 456288 419632 456300
rect 419684 456288 419690 456340
rect 187234 456220 187240 456272
rect 187292 456260 187298 456272
rect 279510 456260 279516 456272
rect 187292 456232 279516 456260
rect 187292 456220 187298 456232
rect 279510 456220 279516 456232
rect 279568 456220 279574 456272
rect 285858 456220 285864 456272
rect 285916 456260 285922 456272
rect 286134 456260 286140 456272
rect 285916 456232 286140 456260
rect 285916 456220 285922 456232
rect 286134 456220 286140 456232
rect 286192 456260 286198 456272
rect 286594 456260 286600 456272
rect 286192 456232 286600 456260
rect 286192 456220 286198 456232
rect 286594 456220 286600 456232
rect 286652 456220 286658 456272
rect 287054 456220 287060 456272
rect 287112 456260 287118 456272
rect 287974 456260 287980 456272
rect 287112 456232 287980 456260
rect 287112 456220 287118 456232
rect 287974 456220 287980 456232
rect 288032 456220 288038 456272
rect 288434 456220 288440 456272
rect 288492 456260 288498 456272
rect 289446 456260 289452 456272
rect 288492 456232 289452 456260
rect 288492 456220 288498 456232
rect 289446 456220 289452 456232
rect 289504 456220 289510 456272
rect 303614 456220 303620 456272
rect 303672 456260 303678 456272
rect 304258 456260 304264 456272
rect 303672 456232 304264 456260
rect 303672 456220 303678 456232
rect 304258 456220 304264 456232
rect 304316 456220 304322 456272
rect 304994 456220 305000 456272
rect 305052 456260 305058 456272
rect 305638 456260 305644 456272
rect 305052 456232 305644 456260
rect 305052 456220 305058 456232
rect 305638 456220 305644 456232
rect 305696 456220 305702 456272
rect 310606 456220 310612 456272
rect 310664 456260 310670 456272
rect 311158 456260 311164 456272
rect 310664 456232 311164 456260
rect 310664 456220 310670 456232
rect 311158 456220 311164 456232
rect 311216 456220 311222 456272
rect 317322 456220 317328 456272
rect 317380 456260 317386 456272
rect 323210 456260 323216 456272
rect 317380 456232 323216 456260
rect 317380 456220 317386 456232
rect 323210 456220 323216 456232
rect 323268 456220 323274 456272
rect 419534 456220 419540 456272
rect 419592 456260 419598 456272
rect 437474 456260 437480 456272
rect 419592 456232 437480 456260
rect 419592 456220 419598 456232
rect 437474 456220 437480 456232
rect 437532 456220 437538 456272
rect 162118 456152 162124 456204
rect 162176 456192 162182 456204
rect 367830 456192 367836 456204
rect 162176 456164 367836 456192
rect 162176 456152 162182 456164
rect 367830 456152 367836 456164
rect 367888 456152 367894 456204
rect 379514 456152 379520 456204
rect 379572 456192 379578 456204
rect 380342 456192 380348 456204
rect 379572 456164 380348 456192
rect 379572 456152 379578 456164
rect 380342 456152 380348 456164
rect 380400 456152 380406 456204
rect 380894 456152 380900 456204
rect 380952 456192 380958 456204
rect 381814 456192 381820 456204
rect 380952 456164 381820 456192
rect 380952 456152 380958 456164
rect 381814 456152 381820 456164
rect 381872 456152 381878 456204
rect 386138 456152 386144 456204
rect 386196 456192 386202 456204
rect 387058 456192 387064 456204
rect 386196 456164 387064 456192
rect 386196 456152 386202 456164
rect 387058 456152 387064 456164
rect 387116 456152 387122 456204
rect 419718 456192 419724 456204
rect 412606 456164 419724 456192
rect 11790 456084 11796 456136
rect 11848 456124 11854 456136
rect 222194 456124 222200 456136
rect 11848 456096 222200 456124
rect 11848 456084 11854 456096
rect 222194 456084 222200 456096
rect 222252 456084 222258 456136
rect 254026 456084 254032 456136
rect 254084 456124 254090 456136
rect 254486 456124 254492 456136
rect 254084 456096 254492 456124
rect 254084 456084 254090 456096
rect 254486 456084 254492 456096
rect 254544 456084 254550 456136
rect 255406 456084 255412 456136
rect 255464 456124 255470 456136
rect 256326 456124 256332 456136
rect 255464 456096 256332 456124
rect 255464 456084 255470 456096
rect 256326 456084 256332 456096
rect 256384 456084 256390 456136
rect 258166 456084 258172 456136
rect 258224 456124 258230 456136
rect 258534 456124 258540 456136
rect 258224 456096 258540 456124
rect 258224 456084 258230 456096
rect 258534 456084 258540 456096
rect 258592 456084 258598 456136
rect 270678 456084 270684 456136
rect 270736 456124 270742 456136
rect 271414 456124 271420 456136
rect 270736 456096 271420 456124
rect 270736 456084 270742 456096
rect 271414 456084 271420 456096
rect 271472 456084 271478 456136
rect 271874 456084 271880 456136
rect 271932 456124 271938 456136
rect 272518 456124 272524 456136
rect 271932 456096 272524 456124
rect 271932 456084 271938 456096
rect 272518 456084 272524 456096
rect 272576 456084 272582 456136
rect 273254 456084 273260 456136
rect 273312 456124 273318 456136
rect 273990 456124 273996 456136
rect 273312 456096 273996 456124
rect 273312 456084 273318 456096
rect 273990 456084 273996 456096
rect 274048 456084 274054 456136
rect 277394 456084 277400 456136
rect 277452 456124 277458 456136
rect 278406 456124 278412 456136
rect 277452 456096 278412 456124
rect 277452 456084 277458 456096
rect 278406 456084 278412 456096
rect 278464 456084 278470 456136
rect 280154 456084 280160 456136
rect 280212 456124 280218 456136
rect 280614 456124 280620 456136
rect 280212 456096 280620 456124
rect 280212 456084 280218 456096
rect 280614 456084 280620 456096
rect 280672 456084 280678 456136
rect 281718 456084 281724 456136
rect 281776 456124 281782 456136
rect 282454 456124 282460 456136
rect 281776 456096 282460 456124
rect 281776 456084 281782 456096
rect 282454 456084 282460 456096
rect 282512 456084 282518 456136
rect 285674 456084 285680 456136
rect 285732 456124 285738 456136
rect 286502 456124 286508 456136
rect 285732 456096 286508 456124
rect 285732 456084 285738 456096
rect 286502 456084 286508 456096
rect 286560 456084 286566 456136
rect 286594 456084 286600 456136
rect 286652 456124 286658 456136
rect 412606 456124 412634 456164
rect 419718 456152 419724 456164
rect 419776 456192 419782 456204
rect 438854 456192 438860 456204
rect 419776 456164 438860 456192
rect 419776 456152 419782 456164
rect 438854 456152 438860 456164
rect 438912 456152 438918 456204
rect 286652 456096 412634 456124
rect 286652 456084 286658 456096
rect 419626 456084 419632 456136
rect 419684 456124 419690 456136
rect 419902 456124 419908 456136
rect 419684 456096 419908 456124
rect 419684 456084 419690 456096
rect 419902 456084 419908 456096
rect 419960 456124 419966 456136
rect 454678 456124 454684 456136
rect 419960 456096 454684 456124
rect 419960 456084 419966 456096
rect 454678 456084 454684 456096
rect 454736 456084 454742 456136
rect 205634 456016 205640 456068
rect 205692 456056 205698 456068
rect 206278 456056 206284 456068
rect 205692 456028 206284 456056
rect 205692 456016 205698 456028
rect 206278 456016 206284 456028
rect 206336 456016 206342 456068
rect 208486 456016 208492 456068
rect 208544 456056 208550 456068
rect 209222 456056 209228 456068
rect 208544 456028 209228 456056
rect 208544 456016 208550 456028
rect 209222 456016 209228 456028
rect 209280 456016 209286 456068
rect 209314 456016 209320 456068
rect 209372 456056 209378 456068
rect 580166 456056 580172 456068
rect 209372 456028 580172 456056
rect 209372 456016 209378 456028
rect 580166 456016 580172 456028
rect 580224 456016 580230 456068
rect 187142 455948 187148 456000
rect 187200 455988 187206 456000
rect 317322 455988 317328 456000
rect 187200 455960 317328 455988
rect 187200 455948 187206 455960
rect 317322 455948 317328 455960
rect 317380 455948 317386 456000
rect 317414 455948 317420 456000
rect 317472 455988 317478 456000
rect 318150 455988 318156 456000
rect 317472 455960 318156 455988
rect 317472 455948 317478 455960
rect 318150 455948 318156 455960
rect 318208 455948 318214 456000
rect 320174 455948 320180 456000
rect 320232 455988 320238 456000
rect 320726 455988 320732 456000
rect 320232 455960 320732 455988
rect 320232 455948 320238 455960
rect 320726 455948 320732 455960
rect 320784 455948 320790 456000
rect 331214 455948 331220 456000
rect 331272 455988 331278 456000
rect 331766 455988 331772 456000
rect 331272 455960 331772 455988
rect 331272 455948 331278 455960
rect 331766 455948 331772 455960
rect 331824 455948 331830 456000
rect 332594 455948 332600 456000
rect 332652 455988 332658 456000
rect 333238 455988 333244 456000
rect 332652 455960 333244 455988
rect 332652 455948 332658 455960
rect 333238 455948 333244 455960
rect 333296 455948 333302 456000
rect 335354 455948 335360 456000
rect 335412 455988 335418 456000
rect 335814 455988 335820 456000
rect 335412 455960 335820 455988
rect 335412 455948 335418 455960
rect 335814 455948 335820 455960
rect 335872 455948 335878 456000
rect 336734 455948 336740 456000
rect 336792 455988 336798 456000
rect 337286 455988 337292 456000
rect 336792 455960 337292 455988
rect 336792 455948 336798 455960
rect 337286 455948 337292 455960
rect 337344 455948 337350 456000
rect 338114 455948 338120 456000
rect 338172 455988 338178 456000
rect 339126 455988 339132 456000
rect 338172 455960 339132 455988
rect 338172 455948 338178 455960
rect 339126 455948 339132 455960
rect 339184 455948 339190 456000
rect 347774 455948 347780 456000
rect 347832 455988 347838 456000
rect 348694 455988 348700 456000
rect 347832 455960 348700 455988
rect 347832 455948 347838 455960
rect 348694 455948 348700 455960
rect 348752 455948 348758 456000
rect 351914 455948 351920 456000
rect 351972 455988 351978 456000
rect 352374 455988 352380 456000
rect 351972 455960 352380 455988
rect 351972 455948 351978 455960
rect 352374 455948 352380 455960
rect 352432 455948 352438 456000
rect 354674 455948 354680 456000
rect 354732 455988 354738 456000
rect 355318 455988 355324 456000
rect 354732 455960 355324 455988
rect 354732 455948 354738 455960
rect 355318 455948 355324 455960
rect 355376 455948 355382 456000
rect 357434 455948 357440 456000
rect 357492 455988 357498 456000
rect 358262 455988 358268 456000
rect 357492 455960 358268 455988
rect 357492 455948 357498 455960
rect 358262 455948 358268 455960
rect 358320 455948 358326 456000
rect 364334 455948 364340 456000
rect 364392 455988 364398 456000
rect 364886 455988 364892 456000
rect 364392 455960 364892 455988
rect 364392 455948 364398 455960
rect 364886 455948 364892 455960
rect 364944 455948 364950 456000
rect 205818 455880 205824 455932
rect 205876 455920 205882 455932
rect 206646 455920 206652 455932
rect 205876 455892 206652 455920
rect 205876 455880 205882 455892
rect 206646 455880 206652 455892
rect 206704 455880 206710 455932
rect 209866 455880 209872 455932
rect 209924 455920 209930 455932
rect 210694 455920 210700 455932
rect 209924 455892 210700 455920
rect 209924 455880 209930 455892
rect 210694 455880 210700 455892
rect 210752 455880 210758 455932
rect 211246 455880 211252 455932
rect 211304 455920 211310 455932
rect 212166 455920 212172 455932
rect 211304 455892 212172 455920
rect 211304 455880 211310 455892
rect 212166 455880 212172 455892
rect 212224 455880 212230 455932
rect 280798 455880 280804 455932
rect 280856 455920 280862 455932
rect 419534 455920 419540 455932
rect 280856 455892 419540 455920
rect 280856 455880 280862 455892
rect 419534 455880 419540 455892
rect 419592 455920 419598 455932
rect 419810 455920 419816 455932
rect 419592 455892 419816 455920
rect 419592 455880 419598 455892
rect 419810 455880 419816 455892
rect 419868 455880 419874 455932
rect 184474 455812 184480 455864
rect 184532 455852 184538 455864
rect 363138 455852 363144 455864
rect 184532 455824 363144 455852
rect 184532 455812 184538 455824
rect 363138 455812 363144 455824
rect 363196 455812 363202 455864
rect 184382 455744 184388 455796
rect 184440 455784 184446 455796
rect 368934 455784 368940 455796
rect 184440 455756 368940 455784
rect 184440 455744 184446 455756
rect 368934 455744 368940 455756
rect 368992 455744 368998 455796
rect 204714 455676 204720 455728
rect 204772 455716 204778 455728
rect 209314 455716 209320 455728
rect 204772 455688 209320 455716
rect 204772 455676 204778 455688
rect 209314 455676 209320 455688
rect 209372 455676 209378 455728
rect 209406 455676 209412 455728
rect 209464 455716 209470 455728
rect 391290 455716 391296 455728
rect 209464 455688 391296 455716
rect 209464 455676 209470 455688
rect 391290 455676 391296 455688
rect 391348 455676 391354 455728
rect 202506 455608 202512 455660
rect 202564 455648 202570 455660
rect 395430 455648 395436 455660
rect 202564 455620 395436 455648
rect 202564 455608 202570 455620
rect 395430 455608 395436 455620
rect 395488 455608 395494 455660
rect 201770 455540 201776 455592
rect 201828 455580 201834 455592
rect 209406 455580 209412 455592
rect 201828 455552 209412 455580
rect 201828 455540 201834 455552
rect 209406 455540 209412 455552
rect 209464 455540 209470 455592
rect 209498 455540 209504 455592
rect 209556 455580 209562 455592
rect 395338 455580 395344 455592
rect 209556 455552 395344 455580
rect 209556 455540 209562 455552
rect 395338 455540 395344 455552
rect 395396 455540 395402 455592
rect 201034 455472 201040 455524
rect 201092 455512 201098 455524
rect 396718 455512 396724 455524
rect 201092 455484 396724 455512
rect 201092 455472 201098 455484
rect 396718 455472 396724 455484
rect 396776 455472 396782 455524
rect 198458 455404 198464 455456
rect 198516 455444 198522 455456
rect 562318 455444 562324 455456
rect 198516 455416 562324 455444
rect 198516 455404 198522 455416
rect 562318 455404 562324 455416
rect 562376 455404 562382 455456
rect 157978 454996 157984 455048
rect 158036 455036 158042 455048
rect 367462 455036 367468 455048
rect 158036 455008 367468 455036
rect 158036 454996 158042 455008
rect 367462 454996 367468 455008
rect 367520 454996 367526 455048
rect 181346 454928 181352 454980
rect 181404 454968 181410 454980
rect 227990 454968 227996 454980
rect 181404 454940 227996 454968
rect 181404 454928 181410 454940
rect 227990 454928 227996 454940
rect 228048 454928 228054 454980
rect 184014 454860 184020 454912
rect 184072 454900 184078 454912
rect 227254 454900 227260 454912
rect 184072 454872 227260 454900
rect 184072 454860 184078 454872
rect 227254 454860 227260 454872
rect 227312 454860 227318 454912
rect 368750 454860 368756 454912
rect 368808 454900 368814 454912
rect 402514 454900 402520 454912
rect 368808 454872 402520 454900
rect 368808 454860 368814 454872
rect 402514 454860 402520 454872
rect 402572 454860 402578 454912
rect 188706 454792 188712 454844
rect 188764 454832 188770 454844
rect 262582 454832 262588 454844
rect 188764 454804 262588 454832
rect 188764 454792 188770 454804
rect 262582 454792 262588 454804
rect 262640 454792 262646 454844
rect 357894 454792 357900 454844
rect 357952 454832 357958 454844
rect 402790 454832 402796 454844
rect 357952 454804 402796 454832
rect 357952 454792 357958 454804
rect 402790 454792 402796 454804
rect 402848 454792 402854 454844
rect 188798 454724 188804 454776
rect 188856 454764 188862 454776
rect 264054 454764 264060 454776
rect 188856 454736 264060 454764
rect 188856 454724 188862 454736
rect 264054 454724 264060 454736
rect 264112 454724 264118 454776
rect 343174 454724 343180 454776
rect 343232 454764 343238 454776
rect 405090 454764 405096 454776
rect 343232 454736 405096 454764
rect 343232 454724 343238 454736
rect 405090 454724 405096 454736
rect 405148 454724 405154 454776
rect 111702 454656 111708 454708
rect 111760 454696 111766 454708
rect 366358 454696 366364 454708
rect 111760 454668 366364 454696
rect 111760 454656 111766 454668
rect 366358 454656 366364 454668
rect 366416 454656 366422 454708
rect 383286 454656 383292 454708
rect 383344 454696 383350 454708
rect 525794 454696 525800 454708
rect 383344 454668 525800 454696
rect 383344 454656 383350 454668
rect 525794 454656 525800 454668
rect 525852 454656 525858 454708
rect 187510 454588 187516 454640
rect 187568 454628 187574 454640
rect 268102 454628 268108 454640
rect 187568 454600 268108 454628
rect 187568 454588 187574 454600
rect 268102 454588 268108 454600
rect 268160 454588 268166 454640
rect 333606 454588 333612 454640
rect 333664 454628 333670 454640
rect 404998 454628 405004 454640
rect 333664 454600 405004 454628
rect 333664 454588 333670 454600
rect 404998 454588 405004 454600
rect 405056 454588 405062 454640
rect 202874 454520 202880 454572
rect 202932 454560 202938 454572
rect 390278 454560 390284 454572
rect 202932 454532 390284 454560
rect 202932 454520 202938 454532
rect 390278 454520 390284 454532
rect 390336 454520 390342 454572
rect 200298 454452 200304 454504
rect 200356 454492 200362 454504
rect 392670 454492 392676 454504
rect 200356 454464 392676 454492
rect 200356 454452 200362 454464
rect 392670 454452 392676 454464
rect 392728 454452 392734 454504
rect 199194 454384 199200 454436
rect 199252 454424 199258 454436
rect 394050 454424 394056 454436
rect 199252 454396 394056 454424
rect 199252 454384 199258 454396
rect 394050 454384 394056 454396
rect 394108 454384 394114 454436
rect 354950 454316 354956 454368
rect 355008 454356 355014 454368
rect 402698 454356 402704 454368
rect 355008 454328 402704 454356
rect 355008 454316 355014 454328
rect 402698 454316 402704 454328
rect 402756 454316 402762 454368
rect 14458 454248 14464 454300
rect 14516 454288 14522 454300
rect 233878 454288 233884 454300
rect 14516 454260 233884 454288
rect 14516 454248 14522 454260
rect 233878 454248 233884 454260
rect 233936 454248 233942 454300
rect 327258 454248 327264 454300
rect 327316 454288 327322 454300
rect 407758 454288 407764 454300
rect 327316 454260 407764 454288
rect 327316 454248 327322 454260
rect 407758 454248 407764 454260
rect 407816 454248 407822 454300
rect 10318 454180 10324 454232
rect 10376 454220 10382 454232
rect 231302 454220 231308 454232
rect 10376 454192 231308 454220
rect 10376 454180 10382 454192
rect 231302 454180 231308 454192
rect 231360 454180 231366 454232
rect 323946 454180 323952 454232
rect 324004 454220 324010 454232
rect 407942 454220 407948 454232
rect 324004 454192 407948 454220
rect 324004 454180 324010 454192
rect 407942 454180 407948 454192
rect 408000 454180 408006 454232
rect 7558 454112 7564 454164
rect 7616 454152 7622 454164
rect 233510 454152 233516 454164
rect 7616 454124 233516 454152
rect 7616 454112 7622 454124
rect 233510 454112 233516 454124
rect 233568 454112 233574 454164
rect 293770 454112 293776 454164
rect 293828 454152 293834 454164
rect 410518 454152 410524 454164
rect 293828 454124 410524 454152
rect 293828 454112 293834 454124
rect 410518 454112 410524 454124
rect 410576 454112 410582 454164
rect 198090 454044 198096 454096
rect 198148 454084 198154 454096
rect 570598 454084 570604 454096
rect 198148 454056 570604 454084
rect 198148 454044 198154 454056
rect 570598 454044 570604 454056
rect 570656 454044 570662 454096
rect 280522 453636 280528 453688
rect 280580 453676 280586 453688
rect 393958 453676 393964 453688
rect 280580 453648 393964 453676
rect 280580 453636 280586 453648
rect 393958 453636 393964 453648
rect 394016 453636 394022 453688
rect 200850 453568 200856 453620
rect 200908 453608 200914 453620
rect 371050 453608 371056 453620
rect 200908 453580 371056 453608
rect 200908 453568 200914 453580
rect 371050 453568 371056 453580
rect 371108 453568 371114 453620
rect 50982 453500 50988 453552
rect 51040 453540 51046 453552
rect 284570 453540 284576 453552
rect 51040 453512 284576 453540
rect 51040 453500 51046 453512
rect 284570 453500 284576 453512
rect 284628 453500 284634 453552
rect 56502 453432 56508 453484
rect 56560 453472 56566 453484
rect 293402 453472 293408 453484
rect 56560 453444 293408 453472
rect 56560 453432 56566 453444
rect 293402 453432 293408 453444
rect 293460 453432 293466 453484
rect 361114 453432 361120 453484
rect 361172 453472 361178 453484
rect 402606 453472 402612 453484
rect 361172 453444 402612 453472
rect 361172 453432 361178 453444
rect 402606 453432 402612 453444
rect 402664 453432 402670 453484
rect 59262 453364 59268 453416
rect 59320 453404 59326 453416
rect 297818 453404 297824 453416
rect 59320 453376 297824 453404
rect 59320 453364 59326 453376
rect 297818 453364 297824 453376
rect 297876 453364 297882 453416
rect 362586 453364 362592 453416
rect 362644 453404 362650 453416
rect 410702 453404 410708 453416
rect 362644 453376 410708 453404
rect 362644 453364 362650 453376
rect 410702 453364 410708 453376
rect 410760 453364 410766 453416
rect 62022 453296 62028 453348
rect 62080 453336 62086 453348
rect 301866 453336 301872 453348
rect 62080 453308 301872 453336
rect 62080 453296 62086 453308
rect 301866 453296 301872 453308
rect 301924 453296 301930 453348
rect 346394 453296 346400 453348
rect 346452 453336 346458 453348
rect 405274 453336 405280 453348
rect 346452 453308 405280 453336
rect 346452 453296 346458 453308
rect 405274 453296 405280 453308
rect 405332 453296 405338 453348
rect 337194 453228 337200 453280
rect 337252 453268 337258 453280
rect 405366 453268 405372 453280
rect 337252 453240 405372 453268
rect 337252 453228 337258 453240
rect 405366 453228 405372 453240
rect 405424 453228 405430 453280
rect 193858 453160 193864 453212
rect 193916 453200 193922 453212
rect 224954 453200 224960 453212
rect 193916 453172 224960 453200
rect 193916 453160 193922 453172
rect 224954 453160 224960 453172
rect 225012 453160 225018 453212
rect 324314 453160 324320 453212
rect 324372 453200 324378 453212
rect 324682 453200 324688 453212
rect 324372 453172 324688 453200
rect 324372 453160 324378 453172
rect 324682 453160 324688 453172
rect 324740 453160 324746 453212
rect 344922 453160 344928 453212
rect 344980 453200 344986 453212
rect 413370 453200 413376 453212
rect 344980 453172 413376 453200
rect 344980 453160 344986 453172
rect 413370 453160 413376 453172
rect 413428 453160 413434 453212
rect 191006 453092 191012 453144
rect 191064 453132 191070 453144
rect 229738 453132 229744 453144
rect 191064 453104 229744 453132
rect 191064 453092 191070 453104
rect 229738 453092 229744 453104
rect 229796 453092 229802 453144
rect 240226 453092 240232 453144
rect 240284 453132 240290 453144
rect 240870 453132 240876 453144
rect 240284 453104 240876 453132
rect 240284 453092 240290 453104
rect 240870 453092 240876 453104
rect 240928 453092 240934 453144
rect 241606 453092 241612 453144
rect 241664 453132 241670 453144
rect 242342 453132 242348 453144
rect 241664 453104 242348 453132
rect 241664 453092 241670 453104
rect 242342 453092 242348 453104
rect 242400 453092 242406 453144
rect 245746 453092 245752 453144
rect 245804 453132 245810 453144
rect 246390 453132 246396 453144
rect 245804 453104 246396 453132
rect 245804 453092 245810 453104
rect 246390 453092 246396 453104
rect 246448 453092 246454 453144
rect 247034 453092 247040 453144
rect 247092 453132 247098 453144
rect 247862 453132 247868 453144
rect 247092 453104 247868 453132
rect 247092 453092 247098 453104
rect 247862 453092 247868 453104
rect 247920 453092 247926 453144
rect 324498 453092 324504 453144
rect 324556 453132 324562 453144
rect 324774 453132 324780 453144
rect 324556 453104 324780 453132
rect 324556 453092 324562 453104
rect 324774 453092 324780 453104
rect 324832 453092 324838 453144
rect 330570 453092 330576 453144
rect 330628 453132 330634 453144
rect 405182 453132 405188 453144
rect 330628 453104 405188 453132
rect 330628 453092 330634 453104
rect 405182 453092 405188 453104
rect 405240 453092 405246 453144
rect 185394 453024 185400 453076
rect 185452 453064 185458 453076
rect 229370 453064 229376 453076
rect 185452 453036 229376 453064
rect 185452 453024 185458 453036
rect 229370 453024 229376 453036
rect 229428 453024 229434 453076
rect 237466 453024 237472 453076
rect 237524 453064 237530 453076
rect 238294 453064 238300 453076
rect 237524 453036 238300 453064
rect 237524 453024 237530 453036
rect 238294 453024 238300 453036
rect 238352 453024 238358 453076
rect 238754 453024 238760 453076
rect 238812 453064 238818 453076
rect 239398 453064 239404 453076
rect 238812 453036 239404 453064
rect 238812 453024 238818 453036
rect 239398 453024 239404 453036
rect 239456 453024 239462 453076
rect 240134 453024 240140 453076
rect 240192 453064 240198 453076
rect 240594 453064 240600 453076
rect 240192 453036 240600 453064
rect 240192 453024 240198 453036
rect 240594 453024 240600 453036
rect 240652 453024 240658 453076
rect 241698 453024 241704 453076
rect 241756 453064 241762 453076
rect 241974 453064 241980 453076
rect 241756 453036 241980 453064
rect 241756 453024 241762 453036
rect 241974 453024 241980 453036
rect 242032 453024 242038 453076
rect 243078 453024 243084 453076
rect 243136 453064 243142 453076
rect 243814 453064 243820 453076
rect 243136 453036 243820 453064
rect 243136 453024 243142 453036
rect 243814 453024 243820 453036
rect 243872 453024 243878 453076
rect 244274 453024 244280 453076
rect 244332 453064 244338 453076
rect 244918 453064 244924 453076
rect 244332 453036 244924 453064
rect 244332 453024 244338 453036
rect 244918 453024 244924 453036
rect 244976 453024 244982 453076
rect 245654 453024 245660 453076
rect 245712 453064 245718 453076
rect 246114 453064 246120 453076
rect 245712 453036 246120 453064
rect 245712 453024 245718 453036
rect 246114 453024 246120 453036
rect 246172 453024 246178 453076
rect 247218 453024 247224 453076
rect 247276 453064 247282 453076
rect 247494 453064 247500 453076
rect 247276 453036 247500 453064
rect 247276 453024 247282 453036
rect 247494 453024 247500 453036
rect 247552 453024 247558 453076
rect 249978 453024 249984 453076
rect 250036 453064 250042 453076
rect 250806 453064 250812 453076
rect 250036 453036 250812 453064
rect 250036 453024 250042 453036
rect 250806 453024 250812 453036
rect 250864 453024 250870 453076
rect 252738 453024 252744 453076
rect 252796 453064 252802 453076
rect 253382 453064 253388 453076
rect 252796 453036 253388 453064
rect 252796 453024 252802 453036
rect 253382 453024 253388 453036
rect 253440 453024 253446 453076
rect 295426 453024 295432 453076
rect 295484 453064 295490 453076
rect 295794 453064 295800 453076
rect 295484 453036 295800 453064
rect 295484 453024 295490 453036
rect 295794 453024 295800 453036
rect 295852 453024 295858 453076
rect 315850 453024 315856 453076
rect 315908 453064 315914 453076
rect 407850 453064 407856 453076
rect 315908 453036 407856 453064
rect 315908 453024 315914 453036
rect 407850 453024 407856 453036
rect 407908 453024 407914 453076
rect 188430 452956 188436 453008
rect 188488 452996 188494 453008
rect 262122 452996 262128 453008
rect 188488 452968 262128 452996
rect 188488 452956 188494 452968
rect 262122 452956 262128 452968
rect 262180 452956 262186 453008
rect 295334 452956 295340 453008
rect 295392 452996 295398 453008
rect 296070 452996 296076 453008
rect 295392 452968 296076 452996
rect 295392 452956 295398 452968
rect 296070 452956 296076 452968
rect 296128 452956 296134 453008
rect 321554 452956 321560 453008
rect 321612 452996 321618 453008
rect 322566 452996 322572 453008
rect 321612 452968 322572 452996
rect 321612 452956 321618 452968
rect 322566 452956 322572 452968
rect 322624 452956 322630 453008
rect 324406 452956 324412 453008
rect 324464 452996 324470 453008
rect 325142 452996 325148 453008
rect 324464 452968 325148 452996
rect 324464 452956 324470 452968
rect 325142 452956 325148 452968
rect 325200 452956 325206 453008
rect 325786 452956 325792 453008
rect 325844 452996 325850 453008
rect 326614 452996 326620 453008
rect 325844 452968 326620 452996
rect 325844 452956 325850 452968
rect 326614 452956 326620 452968
rect 326672 452956 326678 453008
rect 328454 452956 328460 453008
rect 328512 452996 328518 453008
rect 329190 452996 329196 453008
rect 328512 452968 329196 452996
rect 328512 452956 328518 452968
rect 329190 452956 329196 452968
rect 329248 452956 329254 453008
rect 329834 452956 329840 453008
rect 329892 452996 329898 453008
rect 330662 452996 330668 453008
rect 329892 452968 330668 452996
rect 329892 452956 329898 452968
rect 330662 452956 330668 452968
rect 330720 452956 330726 453008
rect 330754 452956 330760 453008
rect 330812 452996 330818 453008
rect 418798 452996 418804 453008
rect 330812 452968 418804 452996
rect 330812 452956 330818 452968
rect 418798 452956 418804 452968
rect 418856 452956 418862 453008
rect 188062 452888 188068 452940
rect 188120 452928 188126 452940
rect 261754 452928 261760 452940
rect 188120 452900 261760 452928
rect 188120 452888 188126 452900
rect 261754 452888 261760 452900
rect 261812 452888 261818 452940
rect 291930 452888 291936 452940
rect 291988 452928 291994 452940
rect 391198 452928 391204 452940
rect 291988 452900 391204 452928
rect 291988 452888 291994 452900
rect 391198 452888 391204 452900
rect 391256 452888 391262 452940
rect 188522 452820 188528 452872
rect 188580 452860 188586 452872
rect 265802 452860 265808 452872
rect 188580 452832 265808 452860
rect 188580 452820 188586 452832
rect 265802 452820 265808 452832
rect 265860 452820 265866 452872
rect 298186 452820 298192 452872
rect 298244 452860 298250 452872
rect 402422 452860 402428 452872
rect 298244 452832 402428 452860
rect 298244 452820 298250 452832
rect 402422 452820 402428 452832
rect 402480 452820 402486 452872
rect 185486 452752 185492 452804
rect 185544 452792 185550 452804
rect 262214 452792 262220 452804
rect 185544 452764 262220 452792
rect 185544 452752 185550 452764
rect 262214 452752 262220 452764
rect 262272 452752 262278 452804
rect 283466 452752 283472 452804
rect 283524 452792 283530 452804
rect 392578 452792 392584 452804
rect 283524 452764 392584 452792
rect 283524 452752 283530 452764
rect 392578 452752 392584 452764
rect 392636 452752 392642 452804
rect 185578 452684 185584 452736
rect 185636 452724 185642 452736
rect 263962 452724 263968 452736
rect 185636 452696 263968 452724
rect 185636 452684 185642 452696
rect 263962 452684 263968 452696
rect 264020 452684 264026 452736
rect 279050 452684 279056 452736
rect 279108 452724 279114 452736
rect 390094 452724 390100 452736
rect 279108 452696 390100 452724
rect 279108 452684 279114 452696
rect 390094 452684 390100 452696
rect 390152 452684 390158 452736
rect 191558 452616 191564 452668
rect 191616 452656 191622 452668
rect 270954 452656 270960 452668
rect 191616 452628 270960 452656
rect 191616 452616 191622 452628
rect 270954 452616 270960 452628
rect 271012 452616 271018 452668
rect 325786 452616 325792 452668
rect 325844 452656 325850 452668
rect 330754 452656 330760 452668
rect 325844 452628 330760 452656
rect 325844 452616 325850 452628
rect 330754 452616 330760 452628
rect 330812 452616 330818 452668
rect 371234 452616 371240 452668
rect 371292 452656 371298 452668
rect 372246 452656 372252 452668
rect 371292 452628 372252 452656
rect 371292 452616 371298 452628
rect 372246 452616 372252 452628
rect 372304 452616 372310 452668
rect 376754 452616 376760 452668
rect 376812 452656 376818 452668
rect 377398 452656 377404 452668
rect 376812 452628 377404 452656
rect 376812 452616 376818 452628
rect 377398 452616 377404 452628
rect 377456 452616 377462 452668
rect 378134 452616 378140 452668
rect 378192 452656 378198 452668
rect 378870 452656 378876 452668
rect 378192 452628 378876 452656
rect 378192 452616 378198 452628
rect 378870 452616 378876 452628
rect 378928 452616 378934 452668
rect 386138 452616 386144 452668
rect 386196 452656 386202 452668
rect 390646 452656 390652 452668
rect 386196 452628 390652 452656
rect 386196 452616 386202 452628
rect 390646 452616 390652 452628
rect 390704 452616 390710 452668
rect 235258 452548 235264 452600
rect 235316 452588 235322 452600
rect 236362 452588 236368 452600
rect 235316 452560 236368 452588
rect 235316 452548 235322 452560
rect 236362 452548 236368 452560
rect 236420 452548 236426 452600
rect 280798 452548 280804 452600
rect 280856 452588 280862 452600
rect 281994 452588 282000 452600
rect 280856 452560 282000 452588
rect 280856 452548 280862 452560
rect 281994 452548 282000 452560
rect 282052 452548 282058 452600
rect 307018 452548 307024 452600
rect 307076 452588 307082 452600
rect 308030 452588 308036 452600
rect 307076 452560 308036 452588
rect 307076 452548 307082 452560
rect 308030 452548 308036 452560
rect 308088 452548 308094 452600
rect 308122 452548 308128 452600
rect 308180 452588 308186 452600
rect 309042 452588 309048 452600
rect 308180 452560 309048 452588
rect 308180 452548 308186 452560
rect 309042 452548 309048 452560
rect 309100 452548 309106 452600
rect 369854 452548 369860 452600
rect 369912 452588 369918 452600
rect 378686 452588 378692 452600
rect 369912 452560 378692 452588
rect 369912 452548 369918 452560
rect 378686 452548 378692 452560
rect 378744 452548 378750 452600
rect 228358 452480 228364 452532
rect 228416 452520 228422 452532
rect 237098 452520 237104 452532
rect 228416 452492 237104 452520
rect 228416 452480 228422 452492
rect 237098 452480 237104 452492
rect 237156 452480 237162 452532
rect 287146 452480 287152 452532
rect 287204 452520 287210 452532
rect 288342 452520 288348 452532
rect 287204 452492 288348 452520
rect 287204 452480 287210 452492
rect 288342 452480 288348 452492
rect 288400 452520 288406 452532
rect 387610 452520 387616 452532
rect 288400 452492 387616 452520
rect 288400 452480 288406 452492
rect 387610 452480 387616 452492
rect 387668 452480 387674 452532
rect 228450 452412 228456 452464
rect 228508 452452 228514 452464
rect 237834 452452 237840 452464
rect 228508 452424 237840 452452
rect 228508 452412 228514 452424
rect 237834 452412 237840 452424
rect 237892 452412 237898 452464
rect 390186 452452 390192 452464
rect 306346 452424 390192 452452
rect 228726 452344 228732 452396
rect 228784 452384 228790 452396
rect 259178 452384 259184 452396
rect 228784 452356 259184 452384
rect 228784 452344 228790 452356
rect 259178 452344 259184 452356
rect 259236 452344 259242 452396
rect 300026 452344 300032 452396
rect 300084 452384 300090 452396
rect 300762 452384 300768 452396
rect 300084 452356 300768 452384
rect 300084 452344 300090 452356
rect 300762 452344 300768 452356
rect 300820 452384 300826 452396
rect 306346 452384 306374 452424
rect 390186 452412 390192 452424
rect 390244 452412 390250 452464
rect 300820 452356 306374 452384
rect 300820 452344 300826 452356
rect 377306 452344 377312 452396
rect 377364 452384 377370 452396
rect 418890 452384 418896 452396
rect 377364 452356 418896 452384
rect 377364 452344 377370 452356
rect 418890 452344 418896 452356
rect 418948 452344 418954 452396
rect 203610 452276 203616 452328
rect 203668 452316 203674 452328
rect 214558 452316 214564 452328
rect 203668 452288 214564 452316
rect 203668 452276 203674 452288
rect 214558 452276 214564 452288
rect 214616 452276 214622 452328
rect 232590 452276 232596 452328
rect 232648 452316 232654 452328
rect 252922 452316 252928 452328
rect 232648 452288 252928 452316
rect 232648 452276 232654 452288
rect 252922 452276 252928 452288
rect 252980 452276 252986 452328
rect 308490 452276 308496 452328
rect 308548 452316 308554 452328
rect 417418 452316 417424 452328
rect 308548 452288 417424 452316
rect 308548 452276 308554 452288
rect 417418 452276 417424 452288
rect 417476 452276 417482 452328
rect 203978 452208 203984 452260
rect 204036 452248 204042 452260
rect 214466 452248 214472 452260
rect 204036 452220 214472 452248
rect 204036 452208 204042 452220
rect 214466 452208 214472 452220
rect 214524 452208 214530 452260
rect 228542 452208 228548 452260
rect 228600 452248 228606 452260
rect 258074 452248 258080 452260
rect 228600 452220 258080 452248
rect 228600 452208 228606 452220
rect 258074 452208 258080 452220
rect 258132 452208 258138 452260
rect 364426 452208 364432 452260
rect 364484 452248 364490 452260
rect 364484 452220 370268 452248
rect 364484 452208 364490 452220
rect 3510 452140 3516 452192
rect 3568 452180 3574 452192
rect 234982 452180 234988 452192
rect 3568 452152 234988 452180
rect 3568 452140 3574 452152
rect 234982 452140 234988 452152
rect 235040 452140 235046 452192
rect 235350 452140 235356 452192
rect 235408 452180 235414 452192
rect 277210 452180 277216 452192
rect 235408 452152 277216 452180
rect 235408 452140 235414 452152
rect 277210 452140 277216 452152
rect 277268 452140 277274 452192
rect 317690 452140 317696 452192
rect 317748 452180 317754 452192
rect 370240 452180 370268 452220
rect 370314 452208 370320 452260
rect 370372 452248 370378 452260
rect 378962 452248 378968 452260
rect 370372 452220 378968 452248
rect 370372 452208 370378 452220
rect 378962 452208 378968 452220
rect 379020 452208 379026 452260
rect 377858 452180 377864 452192
rect 317748 452152 370176 452180
rect 370240 452152 377864 452180
rect 317748 452140 317754 452152
rect 191374 452072 191380 452124
rect 191432 452112 191438 452124
rect 226794 452112 226800 452124
rect 191432 452084 226800 452112
rect 191432 452072 191438 452084
rect 226794 452072 226800 452084
rect 226852 452072 226858 452124
rect 232682 452072 232688 452124
rect 232740 452112 232746 452124
rect 275002 452112 275008 452124
rect 232740 452084 275008 452112
rect 232740 452072 232746 452084
rect 275002 452072 275008 452084
rect 275060 452072 275066 452124
rect 310698 452072 310704 452124
rect 310756 452112 310762 452124
rect 370148 452112 370176 452152
rect 377858 452140 377864 452152
rect 377916 452140 377922 452192
rect 378778 452112 378784 452124
rect 310756 452084 370084 452112
rect 370148 452084 378784 452112
rect 310756 452072 310762 452084
rect 190914 452004 190920 452056
rect 190972 452044 190978 452056
rect 228358 452044 228364 452056
rect 190972 452016 228364 452044
rect 190972 452004 190978 452016
rect 228358 452004 228364 452016
rect 228416 452004 228422 452056
rect 228634 452004 228640 452056
rect 228692 452044 228698 452056
rect 228692 452016 229094 452044
rect 228692 452004 228698 452016
rect 189626 451936 189632 451988
rect 189684 451976 189690 451988
rect 228910 451976 228916 451988
rect 189684 451948 228916 451976
rect 189684 451936 189690 451948
rect 228910 451936 228916 451948
rect 228968 451936 228974 451988
rect 229066 451976 229094 452016
rect 232866 452004 232872 452056
rect 232924 452044 232930 452056
rect 276474 452044 276480 452056
rect 232924 452016 276480 452044
rect 232924 452004 232930 452016
rect 276474 452004 276480 452016
rect 276532 452004 276538 452056
rect 306650 452004 306656 452056
rect 306708 452044 306714 452056
rect 369854 452044 369860 452056
rect 306708 452016 369860 452044
rect 306708 452004 306714 452016
rect 369854 452004 369860 452016
rect 369912 452004 369918 452056
rect 370056 452044 370084 452084
rect 378778 452072 378784 452084
rect 378836 452072 378842 452124
rect 379054 452044 379060 452056
rect 370056 452016 379060 452044
rect 379054 452004 379060 452016
rect 379112 452004 379118 452056
rect 255498 451976 255504 451988
rect 229066 451948 255504 451976
rect 255498 451936 255504 451948
rect 255556 451936 255562 451988
rect 257338 451936 257344 451988
rect 257396 451976 257402 451988
rect 366266 451976 366272 451988
rect 257396 451948 366272 451976
rect 257396 451936 257402 451948
rect 366266 451936 366272 451948
rect 366324 451936 366330 451988
rect 367370 451936 367376 451988
rect 367428 451976 367434 451988
rect 367428 451948 369854 451976
rect 367428 451936 367434 451948
rect 191282 451868 191288 451920
rect 191340 451908 191346 451920
rect 231946 451908 231952 451920
rect 191340 451880 231952 451908
rect 191340 451868 191346 451880
rect 231946 451868 231952 451880
rect 232004 451868 232010 451920
rect 232498 451868 232504 451920
rect 232556 451908 232562 451920
rect 254394 451908 254400 451920
rect 232556 451880 254400 451908
rect 232556 451868 232562 451880
rect 254394 451868 254400 451880
rect 254452 451868 254458 451920
rect 255866 451868 255872 451920
rect 255924 451908 255930 451920
rect 369118 451908 369124 451920
rect 255924 451880 369124 451908
rect 255924 451868 255930 451880
rect 369118 451868 369124 451880
rect 369176 451868 369182 451920
rect 369826 451908 369854 451948
rect 379146 451908 379152 451920
rect 369826 451880 379152 451908
rect 379146 451868 379152 451880
rect 379204 451868 379210 451920
rect 380250 451868 380256 451920
rect 380308 451908 380314 451920
rect 388622 451908 388628 451920
rect 380308 451880 388628 451908
rect 380308 451868 380314 451880
rect 388622 451868 388628 451880
rect 388680 451868 388686 451920
rect 177298 451800 177304 451852
rect 177356 451840 177362 451852
rect 227162 451840 227168 451852
rect 177356 451812 227168 451840
rect 177356 451800 177362 451812
rect 227162 451800 227168 451812
rect 227220 451800 227226 451852
rect 378134 451800 378140 451852
rect 378192 451840 378198 451852
rect 389910 451840 389916 451852
rect 378192 451812 389916 451840
rect 378192 451800 378198 451812
rect 389910 451800 389916 451812
rect 389968 451800 389974 451852
rect 185670 451732 185676 451784
rect 185728 451772 185734 451784
rect 275738 451772 275744 451784
rect 185728 451744 275744 451772
rect 185728 451732 185734 451744
rect 275738 451732 275744 451744
rect 275796 451732 275802 451784
rect 322474 451732 322480 451784
rect 322532 451772 322538 451784
rect 388806 451772 388812 451784
rect 322532 451744 388812 451772
rect 322532 451732 322538 451744
rect 388806 451732 388812 451744
rect 388864 451732 388870 451784
rect 48958 451664 48964 451716
rect 49016 451704 49022 451716
rect 232682 451704 232688 451716
rect 49016 451676 232688 451704
rect 49016 451664 49022 451676
rect 232682 451664 232688 451676
rect 232740 451664 232746 451716
rect 296714 451664 296720 451716
rect 296772 451704 296778 451716
rect 372522 451704 372528 451716
rect 296772 451676 372528 451704
rect 296772 451664 296778 451676
rect 372522 451664 372528 451676
rect 372580 451664 372586 451716
rect 372890 451664 372896 451716
rect 372948 451704 372954 451716
rect 416038 451704 416044 451716
rect 372948 451676 416044 451704
rect 372948 451664 372954 451676
rect 416038 451664 416044 451676
rect 416096 451664 416102 451716
rect 214558 451596 214564 451648
rect 214616 451636 214622 451648
rect 387702 451636 387708 451648
rect 214616 451608 387708 451636
rect 214616 451596 214622 451608
rect 387702 451596 387708 451608
rect 387760 451596 387766 451648
rect 188890 451528 188896 451580
rect 188948 451568 188954 451580
rect 195514 451568 195520 451580
rect 188948 451540 195520 451568
rect 188948 451528 188954 451540
rect 195514 451528 195520 451540
rect 195572 451528 195578 451580
rect 214466 451528 214472 451580
rect 214524 451568 214530 451580
rect 388898 451568 388904 451580
rect 214524 451540 388904 451568
rect 214524 451528 214530 451540
rect 388898 451528 388904 451540
rect 388956 451528 388962 451580
rect 19702 451460 19708 451512
rect 19760 451500 19766 451512
rect 232314 451500 232320 451512
rect 19760 451472 232320 451500
rect 19760 451460 19766 451472
rect 232314 451460 232320 451472
rect 232372 451460 232378 451512
rect 383194 451460 383200 451512
rect 383252 451500 383258 451512
rect 413278 451500 413284 451512
rect 383252 451472 413284 451500
rect 383252 451460 383258 451472
rect 413278 451460 413284 451472
rect 413336 451460 413342 451512
rect 19978 451392 19984 451444
rect 20036 451432 20042 451444
rect 234522 451432 234528 451444
rect 20036 451404 234528 451432
rect 20036 451392 20042 451404
rect 234522 451392 234528 451404
rect 234580 451392 234586 451444
rect 389818 451432 389824 451444
rect 384592 451404 389824 451432
rect 3602 451324 3608 451376
rect 3660 451364 3666 451376
rect 231210 451364 231216 451376
rect 3660 451336 231216 451364
rect 3660 451324 3666 451336
rect 231210 451324 231216 451336
rect 231268 451324 231274 451376
rect 308122 451324 308128 451376
rect 308180 451364 308186 451376
rect 383654 451364 383660 451376
rect 308180 451336 383660 451364
rect 308180 451324 308186 451336
rect 383654 451324 383660 451336
rect 383712 451324 383718 451376
rect 188614 451256 188620 451308
rect 188672 451296 188678 451308
rect 188890 451296 188896 451308
rect 188672 451268 188896 451296
rect 188672 451256 188678 451268
rect 188890 451256 188896 451268
rect 188948 451256 188954 451308
rect 205910 451256 205916 451308
rect 205968 451296 205974 451308
rect 206094 451296 206100 451308
rect 205968 451268 206100 451296
rect 205968 451256 205974 451268
rect 206094 451256 206100 451268
rect 206152 451256 206158 451308
rect 226426 451296 226432 451308
rect 206388 451268 226432 451296
rect 204254 451188 204260 451240
rect 204312 451228 204318 451240
rect 206388 451228 206416 451268
rect 226426 451256 226432 451268
rect 226484 451256 226490 451308
rect 381722 451256 381728 451308
rect 381780 451296 381786 451308
rect 384592 451296 384620 451404
rect 389818 451392 389824 451404
rect 389876 451392 389882 451444
rect 384666 451324 384672 451376
rect 384724 451364 384730 451376
rect 390002 451364 390008 451376
rect 384724 451336 390008 451364
rect 384724 451324 384730 451336
rect 390002 451324 390008 451336
rect 390060 451324 390066 451376
rect 381780 451268 384620 451296
rect 381780 451256 381786 451268
rect 385402 451256 385408 451308
rect 385460 451296 385466 451308
rect 388070 451296 388076 451308
rect 385460 451268 388076 451296
rect 385460 451256 385466 451268
rect 388070 451256 388076 451268
rect 388128 451256 388134 451308
rect 204312 451200 206416 451228
rect 204312 451188 204318 451200
rect 242894 451052 242900 451104
rect 242952 451092 242958 451104
rect 243354 451092 243360 451104
rect 242952 451064 243360 451092
rect 242952 451052 242958 451064
rect 243354 451052 243360 451064
rect 243412 451052 243418 451104
rect 219618 450984 219624 451036
rect 219676 451024 219682 451036
rect 219802 451024 219808 451036
rect 219676 450996 219808 451024
rect 219676 450984 219682 450996
rect 219802 450984 219808 450996
rect 219860 450984 219866 451036
rect 158070 450916 158076 450968
rect 158128 450956 158134 450968
rect 345658 450956 345664 450968
rect 158128 450928 345664 450956
rect 158128 450916 158134 450928
rect 345658 450916 345664 450928
rect 345716 450916 345722 450968
rect 156598 450848 156604 450900
rect 156656 450888 156662 450900
rect 339770 450888 339776 450900
rect 156656 450860 339776 450888
rect 156656 450848 156662 450860
rect 339770 450848 339776 450860
rect 339828 450848 339834 450900
rect 341978 450848 341984 450900
rect 342036 450888 342042 450900
rect 416314 450888 416320 450900
rect 342036 450860 416320 450888
rect 342036 450848 342042 450860
rect 416314 450848 416320 450860
rect 416372 450848 416378 450900
rect 156690 450780 156696 450832
rect 156748 450820 156754 450832
rect 351546 450820 351552 450832
rect 156748 450792 351552 450820
rect 156748 450780 156754 450792
rect 351546 450780 351552 450792
rect 351604 450780 351610 450832
rect 191098 450712 191104 450764
rect 191156 450752 191162 450764
rect 226058 450752 226064 450764
rect 191156 450724 226064 450752
rect 191156 450712 191162 450724
rect 226058 450712 226064 450724
rect 226116 450712 226122 450764
rect 374362 450712 374368 450764
rect 374420 450752 374426 450764
rect 411070 450752 411076 450764
rect 374420 450724 411076 450752
rect 374420 450712 374426 450724
rect 411070 450712 411076 450724
rect 411128 450712 411134 450764
rect 188246 450644 188252 450696
rect 188304 450684 188310 450696
rect 227898 450684 227904 450696
rect 188304 450656 227904 450684
rect 188304 450644 188310 450656
rect 227898 450644 227904 450656
rect 227956 450644 227962 450696
rect 371418 450644 371424 450696
rect 371476 450684 371482 450696
rect 410978 450684 410984 450696
rect 371476 450656 410984 450684
rect 371476 450644 371482 450656
rect 410978 450644 410984 450656
rect 411036 450644 411042 450696
rect 182818 450576 182824 450628
rect 182876 450616 182882 450628
rect 230842 450616 230848 450628
rect 182876 450588 230848 450616
rect 182876 450576 182882 450588
rect 230842 450576 230848 450588
rect 230900 450576 230906 450628
rect 368474 450576 368480 450628
rect 368532 450616 368538 450628
rect 410886 450616 410892 450628
rect 368532 450588 410892 450616
rect 368532 450576 368538 450588
rect 410886 450576 410892 450588
rect 410944 450576 410950 450628
rect 3694 450508 3700 450560
rect 3752 450548 3758 450560
rect 204254 450548 204260 450560
rect 3752 450520 204260 450548
rect 3752 450508 3758 450520
rect 204254 450508 204260 450520
rect 204312 450508 204318 450560
rect 219434 450508 219440 450560
rect 219492 450548 219498 450560
rect 219894 450548 219900 450560
rect 219492 450520 219900 450548
rect 219492 450508 219498 450520
rect 219894 450508 219900 450520
rect 219952 450508 219958 450560
rect 220906 450508 220912 450560
rect 220964 450548 220970 450560
rect 221366 450548 221372 450560
rect 220964 450520 221372 450548
rect 220964 450508 220970 450520
rect 221366 450508 221372 450520
rect 221424 450508 221430 450560
rect 356698 450508 356704 450560
rect 356756 450548 356762 450560
rect 356756 450520 359228 450548
rect 356756 450508 356762 450520
rect 189810 450440 189816 450492
rect 189868 450480 189874 450492
rect 269850 450480 269856 450492
rect 189868 450452 269856 450480
rect 189868 450440 189874 450452
rect 269850 450440 269856 450452
rect 269908 450440 269914 450492
rect 358906 450440 358912 450492
rect 358964 450480 358970 450492
rect 359090 450480 359096 450492
rect 358964 450452 359096 450480
rect 358964 450440 358970 450452
rect 359090 450440 359096 450452
rect 359148 450440 359154 450492
rect 359200 450480 359228 450520
rect 359642 450508 359648 450560
rect 359700 450548 359706 450560
rect 410794 450548 410800 450560
rect 359700 450520 410800 450548
rect 359700 450508 359706 450520
rect 410794 450508 410800 450520
rect 410852 450508 410858 450560
rect 413462 450480 413468 450492
rect 359200 450452 413468 450480
rect 413462 450440 413468 450452
rect 413520 450440 413526 450492
rect 187418 450372 187424 450424
rect 187476 450412 187482 450424
rect 269482 450412 269488 450424
rect 187476 450384 269488 450412
rect 187476 450372 187482 450384
rect 269482 450372 269488 450384
rect 269540 450372 269546 450424
rect 276106 450372 276112 450424
rect 276164 450412 276170 450424
rect 276566 450412 276572 450424
rect 276164 450384 276572 450412
rect 276164 450372 276170 450384
rect 276566 450372 276572 450384
rect 276624 450372 276630 450424
rect 285766 450372 285772 450424
rect 285824 450412 285830 450424
rect 286042 450412 286048 450424
rect 285824 450384 286048 450412
rect 285824 450372 285830 450384
rect 286042 450372 286048 450384
rect 286100 450372 286106 450424
rect 353754 450372 353760 450424
rect 353812 450412 353818 450424
rect 413554 450412 413560 450424
rect 353812 450384 413560 450412
rect 353812 450372 353818 450384
rect 413554 450372 413560 450384
rect 413612 450372 413618 450424
rect 184106 450304 184112 450356
rect 184164 450344 184170 450356
rect 288618 450344 288624 450356
rect 184164 450316 288624 450344
rect 184164 450304 184170 450316
rect 288618 450304 288624 450316
rect 288676 450304 288682 450356
rect 302234 450304 302240 450356
rect 302292 450344 302298 450356
rect 302602 450344 302608 450356
rect 302292 450316 302608 450344
rect 302292 450304 302298 450316
rect 302602 450304 302608 450316
rect 302660 450304 302666 450356
rect 350810 450304 350816 450356
rect 350868 450344 350874 450356
rect 413646 450344 413652 450356
rect 350868 450316 413652 450344
rect 350868 450304 350874 450316
rect 413646 450304 413652 450316
rect 413704 450304 413710 450356
rect 191190 450236 191196 450288
rect 191248 450276 191254 450288
rect 305546 450276 305552 450288
rect 191248 450248 305552 450276
rect 191248 450236 191254 450248
rect 305546 450236 305552 450248
rect 305604 450236 305610 450288
rect 347866 450236 347872 450288
rect 347924 450276 347930 450288
rect 413738 450276 413744 450288
rect 347924 450248 413744 450276
rect 347924 450236 347930 450248
rect 413738 450236 413744 450248
rect 413796 450236 413802 450288
rect 182082 450168 182088 450220
rect 182140 450208 182146 450220
rect 297450 450208 297456 450220
rect 182140 450180 297456 450208
rect 182140 450168 182146 450180
rect 297450 450168 297456 450180
rect 297508 450168 297514 450220
rect 329098 450168 329104 450220
rect 329156 450208 329162 450220
rect 418982 450208 418988 450220
rect 329156 450180 418988 450208
rect 329156 450168 329162 450180
rect 418982 450168 418988 450180
rect 419040 450168 419046 450220
rect 212534 450100 212540 450152
rect 212592 450140 212598 450152
rect 212902 450140 212908 450152
rect 212592 450112 212908 450140
rect 212592 450100 212598 450112
rect 212902 450100 212908 450112
rect 212960 450100 212966 450152
rect 215294 450100 215300 450152
rect 215352 450140 215358 450152
rect 216214 450140 216220 450152
rect 215352 450112 216220 450140
rect 215352 450100 215358 450112
rect 216214 450100 216220 450112
rect 216272 450100 216278 450152
rect 216674 450100 216680 450152
rect 216732 450140 216738 450152
rect 217318 450140 217324 450152
rect 216732 450112 217324 450140
rect 216732 450100 216738 450112
rect 217318 450100 217324 450112
rect 217376 450100 217382 450152
rect 218146 450100 218152 450152
rect 218204 450140 218210 450152
rect 218790 450140 218796 450152
rect 218204 450112 218796 450140
rect 218204 450100 218210 450112
rect 218790 450100 218796 450112
rect 218848 450100 218854 450152
rect 219526 450100 219532 450152
rect 219584 450140 219590 450152
rect 220262 450140 220268 450152
rect 219584 450112 220268 450140
rect 219584 450100 219590 450112
rect 220262 450100 220268 450112
rect 220320 450100 220326 450152
rect 220998 450100 221004 450152
rect 221056 450140 221062 450152
rect 221734 450140 221740 450152
rect 221056 450112 221740 450140
rect 221056 450100 221062 450112
rect 221734 450100 221740 450112
rect 221792 450100 221798 450152
rect 222194 450100 222200 450152
rect 222252 450140 222258 450152
rect 223206 450140 223212 450152
rect 222252 450112 223212 450140
rect 222252 450100 222258 450112
rect 223206 450100 223212 450112
rect 223264 450100 223270 450152
rect 259454 450100 259460 450152
rect 259512 450140 259518 450152
rect 260006 450140 260012 450152
rect 259512 450112 260012 450140
rect 259512 450100 259518 450112
rect 260006 450100 260012 450112
rect 260064 450100 260070 450152
rect 332410 450100 332416 450152
rect 332468 450140 332474 450152
rect 416130 450140 416136 450152
rect 332468 450112 416136 450140
rect 332468 450100 332474 450112
rect 416130 450100 416136 450112
rect 416188 450100 416194 450152
rect 212626 450032 212632 450084
rect 212684 450072 212690 450084
rect 213270 450072 213276 450084
rect 212684 450044 213276 450072
rect 212684 450032 212690 450044
rect 213270 450032 213276 450044
rect 213328 450032 213334 450084
rect 216766 450032 216772 450084
rect 216824 450072 216830 450084
rect 217686 450072 217692 450084
rect 216824 450044 217692 450072
rect 216824 450032 216830 450044
rect 217686 450032 217692 450044
rect 217744 450032 217750 450084
rect 220814 450032 220820 450084
rect 220872 450072 220878 450084
rect 221182 450072 221188 450084
rect 220872 450044 221188 450072
rect 220872 450032 220878 450044
rect 221182 450032 221188 450044
rect 221240 450032 221246 450084
rect 335630 450032 335636 450084
rect 335688 450072 335694 450084
rect 416406 450072 416412 450084
rect 335688 450044 416412 450072
rect 335688 450032 335694 450044
rect 416406 450032 416412 450044
rect 416464 450032 416470 450084
rect 158162 449964 158168 450016
rect 158220 450004 158226 450016
rect 336274 450004 336280 450016
rect 158220 449976 336280 450004
rect 158220 449964 158226 449976
rect 336274 449964 336280 449976
rect 336332 449964 336338 450016
rect 338942 449964 338948 450016
rect 339000 450004 339006 450016
rect 416222 450004 416228 450016
rect 339000 449976 416228 450004
rect 339000 449964 339006 449976
rect 416222 449964 416228 449976
rect 416280 449964 416286 450016
rect 191834 449896 191840 449948
rect 191892 449936 191898 449948
rect 225506 449936 225512 449948
rect 191892 449908 225512 449936
rect 191892 449896 191898 449908
rect 225506 449896 225512 449908
rect 225564 449896 225570 449948
rect 314654 449896 314660 449948
rect 314712 449936 314718 449948
rect 314930 449936 314936 449948
rect 314712 449908 314936 449936
rect 314712 449896 314718 449908
rect 314930 449896 314936 449908
rect 314988 449896 314994 449948
rect 365714 449896 365720 449948
rect 365772 449936 365778 449948
rect 388530 449936 388536 449948
rect 365772 449908 388536 449936
rect 365772 449896 365778 449908
rect 388530 449896 388536 449908
rect 388588 449896 388594 449948
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 193858 449868 193864 449880
rect 3384 449840 193864 449868
rect 3384 449828 3390 449840
rect 193858 449828 193864 449840
rect 193916 449828 193922 449880
rect 387702 449760 387708 449812
rect 387760 449800 387766 449812
rect 388990 449800 388996 449812
rect 387760 449772 388996 449800
rect 387760 449760 387766 449772
rect 388990 449760 388996 449772
rect 389048 449760 389054 449812
rect 349614 449692 349620 449744
rect 349672 449732 349678 449744
rect 405550 449732 405556 449744
rect 349672 449704 405556 449732
rect 349672 449692 349678 449704
rect 405550 449692 405556 449704
rect 405608 449692 405614 449744
rect 190178 449624 190184 449676
rect 190236 449664 190242 449676
rect 263502 449664 263508 449676
rect 190236 449636 263508 449664
rect 190236 449624 190242 449636
rect 263502 449624 263508 449636
rect 263560 449624 263566 449676
rect 312814 449624 312820 449676
rect 312872 449664 312878 449676
rect 407666 449664 407672 449676
rect 312872 449636 407672 449664
rect 312872 449624 312878 449636
rect 407666 449624 407672 449636
rect 407724 449624 407730 449676
rect 189902 449556 189908 449608
rect 189960 449596 189966 449608
rect 267458 449596 267464 449608
rect 189960 449568 267464 449596
rect 189960 449556 189966 449568
rect 267458 449556 267464 449568
rect 267516 449556 267522 449608
rect 268562 449596 268568 449608
rect 267706 449568 268568 449596
rect 189718 449488 189724 449540
rect 189776 449528 189782 449540
rect 267706 449528 267734 449568
rect 268562 449556 268568 449568
rect 268620 449556 268626 449608
rect 309042 449556 309048 449608
rect 309100 449596 309106 449608
rect 408218 449596 408224 449608
rect 309100 449568 408224 449596
rect 309100 449556 309106 449568
rect 408218 449556 408224 449568
rect 408276 449556 408282 449608
rect 189776 449500 267734 449528
rect 189776 449488 189782 449500
rect 388990 449488 388996 449540
rect 389048 449528 389054 449540
rect 580902 449528 580908 449540
rect 389048 449500 580908 449528
rect 389048 449488 389054 449500
rect 580902 449488 580908 449500
rect 580960 449488 580966 449540
rect 188430 447924 188436 447976
rect 188488 447964 188494 447976
rect 188614 447964 188620 447976
rect 188488 447936 188620 447964
rect 188488 447924 188494 447936
rect 188614 447924 188620 447936
rect 188672 447924 188678 447976
rect 188062 446428 188068 446480
rect 188120 446468 188126 446480
rect 188430 446468 188436 446480
rect 188120 446440 188436 446468
rect 188120 446428 188126 446440
rect 188430 446428 188436 446440
rect 188488 446428 188494 446480
rect 388898 442212 388904 442264
rect 388956 442252 388962 442264
rect 580810 442252 580816 442264
rect 388956 442224 580816 442252
rect 388956 442212 388962 442224
rect 580810 442212 580816 442224
rect 580868 442212 580874 442264
rect 390370 422900 390376 422952
rect 390428 422940 390434 422952
rect 580810 422940 580816 422952
rect 390428 422912 580816 422940
rect 390428 422900 390434 422912
rect 580810 422900 580816 422912
rect 580868 422900 580874 422952
rect 394142 419432 394148 419484
rect 394200 419472 394206 419484
rect 580166 419472 580172 419484
rect 394200 419444 580172 419472
rect 394200 419432 394206 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 190822 398800 190828 398812
rect 3384 398772 190828 398800
rect 3384 398760 3390 398772
rect 190822 398760 190828 398772
rect 190880 398760 190886 398812
rect 189534 397400 189540 397452
rect 189592 397440 189598 397452
rect 190822 397440 190828 397452
rect 189592 397412 190828 397440
rect 189592 397400 189598 397412
rect 190822 397400 190828 397412
rect 190880 397400 190886 397452
rect 390278 379448 390284 379500
rect 390336 379488 390342 379500
rect 580166 379488 580172 379500
rect 390336 379460 580172 379488
rect 390336 379448 390342 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3050 372512 3056 372564
rect 3108 372552 3114 372564
rect 190822 372552 190828 372564
rect 3108 372524 190828 372552
rect 3108 372512 3114 372524
rect 190822 372512 190828 372524
rect 190880 372512 190886 372564
rect 399754 365644 399760 365696
rect 399812 365684 399818 365696
rect 580166 365684 580172 365696
rect 399812 365656 580172 365684
rect 399812 365644 399818 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 184014 358748 184020 358760
rect 3384 358720 184020 358748
rect 3384 358708 3390 358720
rect 184014 358708 184020 358720
rect 184072 358708 184078 358760
rect 395430 353200 395436 353252
rect 395488 353240 395494 353252
rect 580166 353240 580172 353252
rect 395488 353212 580172 353240
rect 395488 353200 395494 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 177298 346372 177304 346384
rect 3384 346344 177304 346372
rect 3384 346332 3390 346344
rect 177298 346332 177304 346344
rect 177356 346332 177362 346384
rect 391290 325592 391296 325644
rect 391348 325632 391354 325644
rect 580166 325632 580172 325644
rect 391348 325604 580172 325632
rect 391348 325592 391354 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 2958 320084 2964 320136
rect 3016 320124 3022 320136
rect 188246 320124 188252 320136
rect 3016 320096 188252 320124
rect 3016 320084 3022 320096
rect 188246 320084 188252 320096
rect 188304 320084 188310 320136
rect 403618 313216 403624 313268
rect 403676 313256 403682 313268
rect 580166 313256 580172 313268
rect 403676 313228 580172 313256
rect 403676 313216 403682 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 190914 306320 190920 306332
rect 3384 306292 190920 306320
rect 3384 306280 3390 306292
rect 190914 306280 190920 306292
rect 190972 306280 190978 306332
rect 2866 293904 2872 293956
rect 2924 293944 2930 293956
rect 181346 293944 181352 293956
rect 2924 293916 181352 293944
rect 2924 293904 2930 293916
rect 181346 293904 181352 293916
rect 181404 293904 181410 293956
rect 395338 273164 395344 273216
rect 395396 273204 395402 273216
rect 580166 273204 580172 273216
rect 395396 273176 580172 273204
rect 395396 273164 395402 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 189626 267696 189632 267708
rect 3292 267668 189632 267696
rect 3292 267656 3298 267668
rect 189626 267656 189632 267668
rect 189684 267656 189690 267708
rect 396718 259360 396724 259412
rect 396776 259400 396782 259412
rect 579798 259400 579804 259412
rect 396776 259372 579804 259400
rect 396776 259360 396782 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 3326 255212 3332 255264
rect 3384 255252 3390 255264
rect 190914 255252 190920 255264
rect 3384 255224 190920 255252
rect 3384 255212 3390 255224
rect 190914 255212 190920 255224
rect 190972 255212 190978 255264
rect 186866 250452 186872 250504
rect 186924 250492 186930 250504
rect 218698 250492 218704 250504
rect 186924 250464 218704 250492
rect 186924 250452 186930 250464
rect 218698 250452 218704 250464
rect 218756 250452 218762 250504
rect 378226 249704 378232 249756
rect 378284 249744 378290 249756
rect 386414 249744 386420 249756
rect 378284 249716 386420 249744
rect 378284 249704 378290 249716
rect 386414 249704 386420 249716
rect 386472 249704 386478 249756
rect 386414 248412 386420 248464
rect 386472 248452 386478 248464
rect 389358 248452 389364 248464
rect 386472 248424 389364 248452
rect 386472 248412 386478 248424
rect 389358 248412 389364 248424
rect 389416 248412 389422 248464
rect 216398 248344 216404 248396
rect 216456 248384 216462 248396
rect 236086 248384 236092 248396
rect 216456 248356 236092 248384
rect 216456 248344 216462 248356
rect 236086 248344 236092 248356
rect 236144 248344 236150 248396
rect 313366 248344 313372 248396
rect 313424 248384 313430 248396
rect 358354 248384 358360 248396
rect 313424 248356 358360 248384
rect 313424 248344 313430 248356
rect 358354 248344 358360 248356
rect 358412 248344 358418 248396
rect 383746 248344 383752 248396
rect 383804 248384 383810 248396
rect 389174 248384 389180 248396
rect 383804 248356 389180 248384
rect 383804 248344 383810 248356
rect 389174 248344 389180 248356
rect 389232 248344 389238 248396
rect 217594 248276 217600 248328
rect 217652 248316 217658 248328
rect 237466 248316 237472 248328
rect 217652 248288 237472 248316
rect 217652 248276 217658 248288
rect 237466 248276 237472 248288
rect 237524 248276 237530 248328
rect 314746 248276 314752 248328
rect 314804 248316 314810 248328
rect 360930 248316 360936 248328
rect 314804 248288 360936 248316
rect 314804 248276 314810 248288
rect 360930 248276 360936 248288
rect 360988 248276 360994 248328
rect 385126 248276 385132 248328
rect 385184 248316 385190 248328
rect 389266 248316 389272 248328
rect 385184 248288 389272 248316
rect 385184 248276 385190 248288
rect 389266 248276 389272 248288
rect 389324 248276 389330 248328
rect 217502 248208 217508 248260
rect 217560 248248 217566 248260
rect 238846 248248 238852 248260
rect 217560 248220 238852 248248
rect 217560 248208 217566 248220
rect 238846 248208 238852 248220
rect 238904 248208 238910 248260
rect 316126 248208 316132 248260
rect 316184 248248 316190 248260
rect 363598 248248 363604 248260
rect 316184 248220 363604 248248
rect 316184 248208 316190 248220
rect 363598 248208 363604 248220
rect 363656 248208 363662 248260
rect 382366 248208 382372 248260
rect 382424 248248 382430 248260
rect 388162 248248 388168 248260
rect 382424 248220 388168 248248
rect 382424 248208 382430 248220
rect 388162 248208 388168 248220
rect 388220 248208 388226 248260
rect 217962 248140 217968 248192
rect 218020 248180 218026 248192
rect 240226 248180 240232 248192
rect 218020 248152 240232 248180
rect 218020 248140 218026 248152
rect 240226 248140 240232 248152
rect 240284 248140 240290 248192
rect 311986 248140 311992 248192
rect 312044 248180 312050 248192
rect 359550 248180 359556 248192
rect 312044 248152 359556 248180
rect 312044 248140 312050 248152
rect 359550 248140 359556 248152
rect 359608 248140 359614 248192
rect 379606 248140 379612 248192
rect 379664 248180 379670 248192
rect 391934 248180 391940 248192
rect 379664 248152 391940 248180
rect 379664 248140 379670 248152
rect 391934 248140 391940 248152
rect 391992 248140 391998 248192
rect 182910 248072 182916 248124
rect 182968 248112 182974 248124
rect 201586 248112 201592 248124
rect 182968 248084 201592 248112
rect 182968 248072 182974 248084
rect 201586 248072 201592 248084
rect 201644 248072 201650 248124
rect 217870 248072 217876 248124
rect 217928 248112 217934 248124
rect 241606 248112 241612 248124
rect 217928 248084 241612 248112
rect 217928 248072 217934 248084
rect 241606 248072 241612 248084
rect 241664 248072 241670 248124
rect 276106 248072 276112 248124
rect 276164 248112 276170 248124
rect 357526 248112 357532 248124
rect 276164 248084 357532 248112
rect 276164 248072 276170 248084
rect 357526 248072 357532 248084
rect 357584 248072 357590 248124
rect 380986 248072 380992 248124
rect 381044 248112 381050 248124
rect 390554 248112 390560 248124
rect 381044 248084 390560 248112
rect 381044 248072 381050 248084
rect 390554 248072 390560 248084
rect 390612 248072 390618 248124
rect 181346 248004 181352 248056
rect 181404 248044 181410 248056
rect 200206 248044 200212 248056
rect 181404 248016 200212 248044
rect 181404 248004 181410 248016
rect 200206 248004 200212 248016
rect 200264 248004 200270 248056
rect 217778 248004 217784 248056
rect 217836 248044 217842 248056
rect 242986 248044 242992 248056
rect 217836 248016 242992 248044
rect 217836 248004 217842 248016
rect 242986 248004 242992 248016
rect 243044 248004 243050 248056
rect 305086 248004 305092 248056
rect 305144 248044 305150 248056
rect 402974 248044 402980 248056
rect 305144 248016 402980 248044
rect 305144 248004 305150 248016
rect 402974 248004 402980 248016
rect 403032 248004 403038 248056
rect 179230 247936 179236 247988
rect 179288 247976 179294 247988
rect 204346 247976 204352 247988
rect 179288 247948 204352 247976
rect 179288 247936 179294 247948
rect 204346 247936 204352 247948
rect 204404 247936 204410 247988
rect 219342 247936 219348 247988
rect 219400 247976 219406 247988
rect 245746 247976 245752 247988
rect 219400 247948 245752 247976
rect 219400 247936 219406 247948
rect 245746 247936 245752 247948
rect 245804 247936 245810 247988
rect 299566 247936 299572 247988
rect 299624 247976 299630 247988
rect 304258 247976 304264 247988
rect 299624 247948 304264 247976
rect 299624 247936 299630 247948
rect 304258 247936 304264 247948
rect 304316 247936 304322 247988
rect 306466 247936 306472 247988
rect 306524 247976 306530 247988
rect 407114 247976 407120 247988
rect 306524 247948 407120 247976
rect 306524 247936 306530 247948
rect 407114 247936 407120 247948
rect 407172 247936 407178 247988
rect 174538 247868 174544 247920
rect 174596 247908 174602 247920
rect 207106 247908 207112 247920
rect 174596 247880 207112 247908
rect 174596 247868 174602 247880
rect 207106 247868 207112 247880
rect 207164 247868 207170 247920
rect 217686 247868 217692 247920
rect 217744 247908 217750 247920
rect 244366 247908 244372 247920
rect 217744 247880 244372 247908
rect 217744 247868 217750 247880
rect 244366 247868 244372 247880
rect 244424 247868 244430 247920
rect 307846 247868 307852 247920
rect 307904 247908 307910 247920
rect 409874 247908 409880 247920
rect 307904 247880 409880 247908
rect 307904 247868 307910 247880
rect 409874 247868 409880 247880
rect 409932 247868 409938 247920
rect 175826 247800 175832 247852
rect 175884 247840 175890 247852
rect 208486 247840 208492 247852
rect 175884 247812 208492 247840
rect 175884 247800 175890 247812
rect 208486 247800 208492 247812
rect 208544 247800 208550 247852
rect 216582 247800 216588 247852
rect 216640 247840 216646 247852
rect 248506 247840 248512 247852
rect 216640 247812 248512 247840
rect 216640 247800 216646 247812
rect 248506 247800 248512 247812
rect 248564 247800 248570 247852
rect 309226 247800 309232 247852
rect 309284 247840 309290 247852
rect 414014 247840 414020 247852
rect 309284 247812 414020 247840
rect 309284 247800 309290 247812
rect 414014 247800 414020 247812
rect 414072 247800 414078 247852
rect 1394 247732 1400 247784
rect 1452 247772 1458 247784
rect 193306 247772 193312 247784
rect 1452 247744 193312 247772
rect 1452 247732 1458 247744
rect 193306 247732 193312 247744
rect 193364 247732 193370 247784
rect 215202 247732 215208 247784
rect 215260 247772 215266 247784
rect 247126 247772 247132 247784
rect 215260 247744 247132 247772
rect 215260 247732 215266 247744
rect 247126 247732 247132 247744
rect 247184 247732 247190 247784
rect 267826 247732 267832 247784
rect 267884 247772 267890 247784
rect 356606 247772 356612 247784
rect 267884 247744 356612 247772
rect 267884 247732 267890 247744
rect 356606 247732 356612 247744
rect 356664 247732 356670 247784
rect 387886 247732 387892 247784
rect 387944 247772 387950 247784
rect 558914 247772 558920 247784
rect 387944 247744 558920 247772
rect 387944 247732 387950 247744
rect 558914 247732 558920 247744
rect 558972 247732 558978 247784
rect 14 247664 20 247716
rect 72 247704 78 247716
rect 191926 247704 191932 247716
rect 72 247676 191932 247704
rect 72 247664 78 247676
rect 191926 247664 191932 247676
rect 191984 247664 191990 247716
rect 216490 247664 216496 247716
rect 216548 247704 216554 247716
rect 249886 247704 249892 247716
rect 216548 247676 249892 247704
rect 216548 247664 216554 247676
rect 249886 247664 249892 247676
rect 249944 247664 249950 247716
rect 271966 247664 271972 247716
rect 272024 247704 272030 247716
rect 361666 247704 361672 247716
rect 272024 247676 361672 247704
rect 272024 247664 272030 247676
rect 361666 247664 361672 247676
rect 361724 247664 361730 247716
rect 376846 247664 376852 247716
rect 376904 247704 376910 247716
rect 582374 247704 582380 247716
rect 376904 247676 582380 247704
rect 376904 247664 376910 247676
rect 582374 247664 582380 247676
rect 582432 247664 582438 247716
rect 211246 247596 211252 247648
rect 211304 247636 211310 247648
rect 230566 247636 230572 247648
rect 211304 247608 230572 247636
rect 211304 247596 211310 247608
rect 230566 247596 230572 247608
rect 230624 247596 230630 247648
rect 320266 247596 320272 247648
rect 320324 247636 320330 247648
rect 358170 247636 358176 247648
rect 320324 247608 358176 247636
rect 320324 247596 320330 247608
rect 358170 247596 358176 247608
rect 358228 247596 358234 247648
rect 217410 247528 217416 247580
rect 217468 247568 217474 247580
rect 234706 247568 234712 247580
rect 217468 247540 234712 247568
rect 217468 247528 217474 247540
rect 234706 247528 234712 247540
rect 234764 247528 234770 247580
rect 331306 247528 331312 247580
rect 331364 247568 331370 247580
rect 359458 247568 359464 247580
rect 331364 247540 359464 247568
rect 331364 247528 331370 247540
rect 359458 247528 359464 247540
rect 359516 247528 359522 247580
rect 215294 247460 215300 247512
rect 215352 247500 215358 247512
rect 231946 247500 231952 247512
rect 215352 247472 231952 247500
rect 215352 247460 215358 247472
rect 231946 247460 231952 247472
rect 232004 247460 232010 247512
rect 338206 247460 338212 247512
rect 338264 247500 338270 247512
rect 356698 247500 356704 247512
rect 338264 247472 356704 247500
rect 338264 247460 338270 247472
rect 356698 247460 356704 247472
rect 356756 247460 356762 247512
rect 291286 247120 291292 247172
rect 291344 247160 291350 247172
rect 293218 247160 293224 247172
rect 291344 247132 293224 247160
rect 291344 247120 291350 247132
rect 293218 247120 293224 247132
rect 293276 247120 293282 247172
rect 298186 247120 298192 247172
rect 298244 247160 298250 247172
rect 302878 247160 302884 247172
rect 298244 247132 302884 247160
rect 298244 247120 298250 247132
rect 302878 247120 302884 247132
rect 302936 247120 302942 247172
rect 195238 247052 195244 247104
rect 195296 247092 195302 247104
rect 196066 247092 196072 247104
rect 195296 247064 196072 247092
rect 195296 247052 195302 247064
rect 196066 247052 196072 247064
rect 196124 247052 196130 247104
rect 231118 247052 231124 247104
rect 231176 247092 231182 247104
rect 233326 247092 233332 247104
rect 231176 247064 233332 247092
rect 231176 247052 231182 247064
rect 233326 247052 233332 247064
rect 233384 247052 233390 247104
rect 289906 247052 289912 247104
rect 289964 247092 289970 247104
rect 291838 247092 291844 247104
rect 289964 247064 291844 247092
rect 289964 247052 289970 247064
rect 291838 247052 291844 247064
rect 291896 247052 291902 247104
rect 294046 247052 294052 247104
rect 294104 247092 294110 247104
rect 295978 247092 295984 247104
rect 294104 247064 295984 247092
rect 294104 247052 294110 247064
rect 295978 247052 295984 247064
rect 296036 247052 296042 247104
rect 296806 247052 296812 247104
rect 296864 247092 296870 247104
rect 298738 247092 298744 247104
rect 296864 247064 298744 247092
rect 296864 247052 296870 247064
rect 298738 247052 298744 247064
rect 298796 247052 298802 247104
rect 300946 247052 300952 247104
rect 301004 247092 301010 247104
rect 305638 247092 305644 247104
rect 301004 247064 305644 247092
rect 301004 247052 301010 247064
rect 305638 247052 305644 247064
rect 305696 247052 305702 247104
rect 165614 246304 165620 246356
rect 165672 246344 165678 246356
rect 212626 246344 212632 246356
rect 165672 246316 212632 246344
rect 165672 246304 165678 246316
rect 212626 246304 212632 246316
rect 212684 246304 212690 246356
rect 292666 246304 292672 246356
rect 292724 246344 292730 246356
rect 371234 246344 371240 246356
rect 292724 246316 371240 246344
rect 292724 246304 292730 246316
rect 371234 246304 371240 246316
rect 371292 246304 371298 246356
rect 386414 246304 386420 246356
rect 386472 246344 386478 246356
rect 415394 246344 415400 246356
rect 386472 246316 415400 246344
rect 386472 246304 386478 246316
rect 415394 246304 415400 246316
rect 415452 246304 415458 246356
rect 387058 245624 387064 245676
rect 387116 245664 387122 245676
rect 387886 245664 387892 245676
rect 387116 245636 387892 245664
rect 387116 245624 387122 245636
rect 387886 245624 387892 245636
rect 387944 245624 387950 245676
rect 392670 245556 392676 245608
rect 392728 245596 392734 245608
rect 580166 245596 580172 245608
rect 392728 245568 580172 245596
rect 392728 245556 392734 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 161474 244876 161480 244928
rect 161532 244916 161538 244928
rect 211154 244916 211160 244928
rect 161532 244888 211160 244916
rect 161532 244876 161538 244888
rect 211154 244876 211160 244888
rect 211212 244876 211218 244928
rect 325786 244876 325792 244928
rect 325844 244916 325850 244928
rect 411898 244916 411904 244928
rect 325844 244888 411904 244916
rect 325844 244876 325850 244888
rect 411898 244876 411904 244888
rect 411956 244876 411962 244928
rect 332686 243584 332692 243636
rect 332744 243624 332750 243636
rect 381538 243624 381544 243636
rect 332744 243596 381544 243624
rect 332744 243584 332750 243596
rect 381538 243584 381544 243596
rect 381596 243584 381602 243636
rect 172514 243516 172520 243568
rect 172572 243556 172578 243568
rect 215386 243556 215392 243568
rect 172572 243528 215392 243556
rect 172572 243516 172578 243528
rect 215386 243516 215392 243528
rect 215444 243516 215450 243568
rect 368566 243516 368572 243568
rect 368624 243556 368630 243568
rect 565814 243556 565820 243568
rect 368624 243528 565820 243556
rect 368624 243516 368630 243528
rect 565814 243516 565820 243528
rect 565872 243516 565878 243568
rect 176654 242156 176660 242208
rect 176712 242196 176718 242208
rect 216766 242196 216772 242208
rect 176712 242168 216772 242196
rect 176712 242156 176718 242168
rect 216766 242156 216772 242168
rect 216824 242156 216830 242208
rect 371326 242156 371332 242208
rect 371384 242196 371390 242208
rect 565078 242196 565084 242208
rect 371384 242168 565084 242196
rect 371384 242156 371390 242168
rect 565078 242156 565084 242168
rect 565136 242156 565142 242208
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 185394 241448 185400 241460
rect 3292 241420 185400 241448
rect 3292 241408 3298 241420
rect 185394 241408 185400 241420
rect 185452 241408 185458 241460
rect 295334 239436 295340 239488
rect 295392 239476 295398 239488
rect 378134 239476 378140 239488
rect 295392 239448 378140 239476
rect 295392 239436 295398 239448
rect 378134 239436 378140 239448
rect 378192 239436 378198 239488
rect 179414 239368 179420 239420
rect 179472 239408 179478 239420
rect 218054 239408 218060 239420
rect 179472 239380 218060 239408
rect 179472 239368 179478 239380
rect 218054 239368 218060 239380
rect 218112 239368 218118 239420
rect 372614 239368 372620 239420
rect 372672 239408 372678 239420
rect 569218 239408 569224 239420
rect 372672 239380 569224 239408
rect 372672 239368 372678 239380
rect 569218 239368 569224 239380
rect 569276 239368 569282 239420
rect 293218 236648 293224 236700
rect 293276 236688 293282 236700
rect 367186 236688 367192 236700
rect 293276 236660 367192 236688
rect 293276 236648 293282 236660
rect 367186 236648 367192 236660
rect 367244 236648 367250 236700
rect 373994 236648 374000 236700
rect 374052 236688 374058 236700
rect 578878 236688 578884 236700
rect 374052 236660 578884 236688
rect 374052 236648 374058 236660
rect 578878 236648 578884 236660
rect 578936 236648 578942 236700
rect 328454 233860 328460 233912
rect 328512 233900 328518 233912
rect 408402 233900 408408 233912
rect 328512 233872 408408 233900
rect 328512 233860 328518 233872
rect 408402 233860 408408 233872
rect 408460 233860 408466 233912
rect 298738 232500 298744 232552
rect 298796 232540 298802 232552
rect 382274 232540 382280 232552
rect 298796 232512 382280 232540
rect 298796 232500 298802 232512
rect 382274 232500 382280 232512
rect 382332 232500 382338 232552
rect 302878 229712 302884 229764
rect 302936 229752 302942 229764
rect 385034 229752 385040 229764
rect 302936 229724 385040 229752
rect 302936 229712 302942 229724
rect 385034 229712 385040 229724
rect 385092 229712 385098 229764
rect 3786 217268 3792 217320
rect 3844 217308 3850 217320
rect 191282 217308 191288 217320
rect 3844 217280 191288 217308
rect 3844 217268 3850 217280
rect 191282 217268 191288 217280
rect 191340 217268 191346 217320
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 187326 215268 187332 215280
rect 3384 215240 187332 215268
rect 3384 215228 3390 215240
rect 187326 215228 187332 215240
rect 187384 215228 187390 215280
rect 394050 206932 394056 206984
rect 394108 206972 394114 206984
rect 579798 206972 579804 206984
rect 394108 206944 579804 206972
rect 394108 206932 394114 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 3326 202784 3332 202836
rect 3384 202824 3390 202836
rect 182818 202824 182824 202836
rect 3384 202796 182824 202824
rect 3384 202784 3390 202796
rect 182818 202784 182824 202796
rect 182876 202784 182882 202836
rect 375374 199384 375380 199436
rect 375432 199424 375438 199436
rect 562410 199424 562416 199436
rect 375432 199396 562416 199424
rect 375432 199384 375438 199396
rect 562410 199384 562416 199396
rect 562468 199384 562474 199436
rect 369854 197956 369860 198008
rect 369912 197996 369918 198008
rect 569954 197996 569960 198008
rect 369912 197968 569960 197996
rect 369912 197956 369918 197968
rect 569954 197956 569960 197968
rect 570012 197956 570018 198008
rect 150986 195984 150992 196036
rect 151044 196024 151050 196036
rect 157334 196024 157340 196036
rect 151044 195996 157340 196024
rect 151044 195984 151050 195996
rect 157334 195984 157340 195996
rect 157392 195984 157398 196036
rect 551002 195984 551008 196036
rect 551060 196024 551066 196036
rect 557534 196024 557540 196036
rect 551060 195996 557540 196024
rect 551060 195984 551066 195996
rect 557534 195984 557540 195996
rect 557592 195984 557598 196036
rect 18414 195508 18420 195560
rect 18472 195548 18478 195560
rect 34514 195548 34520 195560
rect 18472 195520 34520 195548
rect 18472 195508 18478 195520
rect 34514 195508 34520 195520
rect 34572 195508 34578 195560
rect 17126 195440 17132 195492
rect 17184 195480 17190 195492
rect 52454 195480 52460 195492
rect 17184 195452 52460 195480
rect 17184 195440 17190 195452
rect 52454 195440 52460 195452
rect 52512 195440 52518 195492
rect 18690 195372 18696 195424
rect 18748 195412 18754 195424
rect 66254 195412 66260 195424
rect 18748 195384 66260 195412
rect 18748 195372 18754 195384
rect 66254 195372 66260 195384
rect 66312 195372 66318 195424
rect 19610 195304 19616 195356
rect 19668 195344 19674 195356
rect 80146 195344 80152 195356
rect 19668 195316 80152 195344
rect 19668 195304 19674 195316
rect 80146 195304 80152 195316
rect 80204 195304 80210 195356
rect 18506 195236 18512 195288
rect 18564 195276 18570 195288
rect 80054 195276 80060 195288
rect 18564 195248 80060 195276
rect 18564 195236 18570 195248
rect 80054 195236 80060 195248
rect 80112 195236 80118 195288
rect 3694 193808 3700 193860
rect 3752 193848 3758 193860
rect 48958 193848 48964 193860
rect 3752 193820 48964 193848
rect 3752 193808 3758 193820
rect 48958 193808 48964 193820
rect 49016 193808 49022 193860
rect 562318 193128 562324 193180
rect 562376 193168 562382 193180
rect 579614 193168 579620 193180
rect 562376 193140 579620 193168
rect 562376 193128 562382 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 3326 188980 3332 189032
rect 3384 189020 3390 189032
rect 18598 189020 18604 189032
rect 3384 188992 18604 189020
rect 3384 188980 3390 188992
rect 18598 188980 18604 188992
rect 18656 188980 18662 189032
rect 310514 180072 310520 180124
rect 310572 180112 310578 180124
rect 416498 180112 416504 180124
rect 310572 180084 416504 180112
rect 310572 180072 310578 180084
rect 416498 180072 416504 180084
rect 416556 180072 416562 180124
rect 570598 166948 570604 167000
rect 570656 166988 570662 167000
rect 580166 166988 580172 167000
rect 570656 166960 580172 166988
rect 570656 166948 570662 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 573358 153144 573364 153196
rect 573416 153184 573422 153196
rect 580166 153184 580172 153196
rect 573416 153156 580172 153184
rect 573416 153144 573422 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 405642 146888 405648 146940
rect 405700 146928 405706 146940
rect 416774 146928 416780 146940
rect 405700 146900 416780 146928
rect 405700 146888 405706 146900
rect 416774 146888 416780 146900
rect 416832 146888 416838 146940
rect 413922 144848 413928 144900
rect 413980 144888 413986 144900
rect 417142 144888 417148 144900
rect 413980 144860 417148 144888
rect 413980 144848 413986 144860
rect 417142 144848 417148 144860
rect 417200 144848 417206 144900
rect 411162 141380 411168 141432
rect 411220 141420 411226 141432
rect 416774 141420 416780 141432
rect 411220 141392 416780 141420
rect 411220 141380 411226 141392
rect 416774 141380 416780 141392
rect 416832 141380 416838 141432
rect 409782 140020 409788 140072
rect 409840 140060 409846 140072
rect 416774 140060 416780 140072
rect 409840 140032 416780 140060
rect 409840 140020 409846 140032
rect 416774 140020 416780 140032
rect 416832 140020 416838 140072
rect 15930 138252 15936 138304
rect 15988 138292 15994 138304
rect 17862 138292 17868 138304
rect 15988 138264 17868 138292
rect 15988 138252 15994 138264
rect 17862 138252 17868 138264
rect 17920 138252 17926 138304
rect 3050 137912 3056 137964
rect 3108 137952 3114 137964
rect 10318 137952 10324 137964
rect 3108 137924 10324 137952
rect 3108 137912 3114 137924
rect 10318 137912 10324 137924
rect 10376 137912 10382 137964
rect 417142 137300 417148 137352
rect 417200 137340 417206 137352
rect 417602 137340 417608 137352
rect 417200 137312 417608 137340
rect 417200 137300 417206 137312
rect 417602 137300 417608 137312
rect 417660 137300 417666 137352
rect 333974 129004 333980 129056
rect 334032 129044 334038 129056
rect 406378 129044 406384 129056
rect 334032 129016 406384 129044
rect 334032 129004 334038 129016
rect 406378 129004 406384 129016
rect 406436 129004 406442 129056
rect 327074 127576 327080 127628
rect 327132 127616 327138 127628
rect 413830 127616 413836 127628
rect 327132 127588 413836 127616
rect 327132 127576 327138 127588
rect 413830 127576 413836 127588
rect 413888 127576 413894 127628
rect 566458 126896 566464 126948
rect 566516 126936 566522 126948
rect 580166 126936 580172 126948
rect 566516 126908 580172 126936
rect 566516 126896 566522 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 324314 126216 324320 126268
rect 324372 126256 324378 126268
rect 416590 126256 416596 126268
rect 324372 126228 416596 126256
rect 324372 126216 324378 126228
rect 416590 126216 416596 126228
rect 416648 126216 416654 126268
rect 322934 124856 322940 124908
rect 322992 124896 322998 124908
rect 414658 124896 414664 124908
rect 322992 124868 414664 124896
rect 322992 124856 322998 124868
rect 414658 124856 414664 124868
rect 414716 124856 414722 124908
rect 321554 123428 321560 123480
rect 321612 123468 321618 123480
rect 415946 123468 415952 123480
rect 321612 123440 415952 123468
rect 321612 123428 321618 123440
rect 415946 123428 415952 123440
rect 416004 123428 416010 123480
rect 291838 122068 291844 122120
rect 291896 122108 291902 122120
rect 364426 122108 364432 122120
rect 291896 122080 364432 122108
rect 291896 122068 291902 122080
rect 364426 122068 364432 122080
rect 364484 122068 364490 122120
rect 287054 120708 287060 120760
rect 287112 120748 287118 120760
rect 357618 120748 357624 120760
rect 287112 120720 357624 120748
rect 287112 120708 287118 120720
rect 357618 120708 357624 120720
rect 357676 120708 357682 120760
rect 417786 120164 417792 120216
rect 417844 120204 417850 120216
rect 419258 120204 419264 120216
rect 417844 120176 419264 120204
rect 417844 120164 417850 120176
rect 419258 120164 419264 120176
rect 419316 120164 419322 120216
rect 351178 117920 351184 117972
rect 351236 117960 351242 117972
rect 415394 117960 415400 117972
rect 351236 117932 415400 117960
rect 351236 117920 351242 117932
rect 415394 117920 415400 117932
rect 415452 117960 415458 117972
rect 417786 117960 417792 117972
rect 415452 117932 417792 117960
rect 415452 117920 415458 117932
rect 417786 117920 417792 117932
rect 417844 117920 417850 117972
rect 305638 115200 305644 115252
rect 305696 115240 305702 115252
rect 391934 115240 391940 115252
rect 305696 115212 391940 115240
rect 305696 115200 305702 115212
rect 391934 115200 391940 115212
rect 391992 115200 391998 115252
rect 304258 113772 304264 113824
rect 304316 113812 304322 113824
rect 389174 113812 389180 113824
rect 304316 113784 389180 113812
rect 304316 113772 304322 113784
rect 389174 113772 389180 113784
rect 389232 113772 389238 113824
rect 571978 113092 571984 113144
rect 572036 113132 572042 113144
rect 579982 113132 579988 113144
rect 572036 113104 579988 113132
rect 572036 113092 572042 113104
rect 579982 113092 579988 113104
rect 580040 113092 580046 113144
rect 295978 112548 295984 112600
rect 296036 112588 296042 112600
rect 373994 112588 374000 112600
rect 296036 112560 374000 112588
rect 296036 112548 296042 112560
rect 373994 112548 374000 112560
rect 374052 112548 374058 112600
rect 303614 112480 303620 112532
rect 303672 112520 303678 112532
rect 398834 112520 398840 112532
rect 303672 112492 398840 112520
rect 303672 112480 303678 112492
rect 398834 112480 398840 112492
rect 398892 112480 398898 112532
rect 318794 112412 318800 112464
rect 318852 112452 318858 112464
rect 419074 112452 419080 112464
rect 318852 112424 419080 112452
rect 318852 112412 318858 112424
rect 419074 112412 419080 112424
rect 419132 112412 419138 112464
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 19702 111772 19708 111784
rect 3384 111744 19708 111772
rect 3384 111732 3390 111744
rect 19702 111732 19708 111744
rect 19760 111732 19766 111784
rect 288434 111188 288440 111240
rect 288492 111228 288498 111240
rect 360286 111228 360292 111240
rect 288492 111200 360292 111228
rect 288492 111188 288498 111200
rect 360286 111188 360292 111200
rect 360344 111188 360350 111240
rect 302234 111120 302240 111172
rect 302292 111160 302298 111172
rect 396074 111160 396080 111172
rect 302292 111132 396080 111160
rect 302292 111120 302298 111132
rect 396074 111120 396080 111132
rect 396132 111120 396138 111172
rect 317414 111052 317420 111104
rect 317472 111092 317478 111104
rect 418522 111092 418528 111104
rect 317472 111064 418528 111092
rect 317472 111052 317478 111064
rect 418522 111052 418528 111064
rect 418580 111052 418586 111104
rect 417970 109692 417976 109744
rect 418028 109732 418034 109744
rect 451274 109732 451280 109744
rect 418028 109704 451280 109732
rect 418028 109692 418034 109704
rect 451274 109692 451280 109704
rect 451332 109732 451338 109744
rect 452470 109732 452476 109744
rect 451332 109704 452476 109732
rect 451332 109692 451338 109704
rect 452470 109692 452476 109704
rect 452528 109692 452534 109744
rect 418982 109624 418988 109676
rect 419040 109664 419046 109676
rect 480898 109664 480904 109676
rect 419040 109636 480904 109664
rect 419040 109624 419046 109636
rect 480898 109624 480904 109636
rect 480956 109624 480962 109676
rect 416130 109556 416136 109608
rect 416188 109596 416194 109608
rect 483474 109596 483480 109608
rect 416188 109568 483480 109596
rect 416188 109556 416194 109568
rect 483474 109556 483480 109568
rect 483532 109556 483538 109608
rect 416406 109488 416412 109540
rect 416464 109528 416470 109540
rect 485958 109528 485964 109540
rect 416464 109500 485964 109528
rect 416464 109488 416470 109500
rect 485958 109488 485964 109500
rect 486016 109488 486022 109540
rect 416222 109420 416228 109472
rect 416280 109460 416286 109472
rect 488258 109460 488264 109472
rect 416280 109432 488264 109460
rect 416280 109420 416286 109432
rect 488258 109420 488264 109432
rect 488316 109420 488322 109472
rect 416314 109352 416320 109404
rect 416372 109392 416378 109404
rect 491018 109392 491024 109404
rect 416372 109364 491024 109392
rect 416372 109352 416378 109364
rect 491018 109352 491024 109364
rect 491076 109352 491082 109404
rect 413370 109284 413376 109336
rect 413428 109324 413434 109336
rect 493410 109324 493416 109336
rect 413428 109296 493416 109324
rect 413428 109284 413434 109296
rect 493410 109284 493416 109296
rect 493468 109284 493474 109336
rect 413738 109216 413744 109268
rect 413796 109256 413802 109268
rect 495894 109256 495900 109268
rect 413796 109228 495900 109256
rect 413796 109216 413802 109228
rect 495894 109216 495900 109228
rect 495952 109216 495958 109268
rect 413646 109148 413652 109200
rect 413704 109188 413710 109200
rect 498470 109188 498476 109200
rect 413704 109160 498476 109188
rect 413704 109148 413710 109160
rect 498470 109148 498476 109160
rect 498528 109148 498534 109200
rect 388806 109080 388812 109132
rect 388864 109120 388870 109132
rect 476114 109120 476120 109132
rect 388864 109092 476120 109120
rect 388864 109080 388870 109092
rect 476114 109080 476120 109092
rect 476172 109080 476178 109132
rect 410702 109012 410708 109064
rect 410760 109052 410766 109064
rect 508498 109052 508504 109064
rect 410760 109024 508504 109052
rect 410760 109012 410766 109024
rect 508498 109012 508504 109024
rect 508556 109012 508562 109064
rect 113450 108944 113456 108996
rect 113508 108984 113514 108996
rect 184382 108984 184388 108996
rect 113508 108956 184388 108984
rect 113508 108944 113514 108956
rect 184382 108944 184388 108956
rect 184440 108944 184446 108996
rect 111058 108876 111064 108928
rect 111116 108916 111122 108928
rect 184290 108916 184296 108928
rect 111116 108888 184296 108916
rect 111116 108876 111122 108888
rect 184290 108876 184296 108888
rect 184348 108876 184354 108928
rect 108574 108808 108580 108860
rect 108632 108848 108638 108860
rect 184474 108848 184480 108860
rect 108632 108820 184480 108848
rect 108632 108808 108638 108820
rect 184474 108808 184480 108820
rect 184532 108808 184538 108860
rect 413554 108808 413560 108860
rect 413612 108848 413618 108860
rect 500954 108848 500960 108860
rect 413612 108820 500960 108848
rect 413612 108808 413618 108820
rect 500954 108808 500960 108820
rect 501012 108808 501018 108860
rect 105998 108740 106004 108792
rect 106056 108780 106062 108792
rect 184198 108780 184204 108792
rect 106056 108752 184204 108780
rect 106056 108740 106062 108752
rect 184198 108740 184204 108752
rect 184256 108740 184262 108792
rect 413462 108740 413468 108792
rect 413520 108780 413526 108792
rect 503438 108780 503444 108792
rect 413520 108752 503444 108780
rect 413520 108740 413526 108752
rect 503438 108740 503444 108752
rect 503496 108740 503502 108792
rect 100938 108672 100944 108724
rect 100996 108712 101002 108724
rect 184658 108712 184664 108724
rect 100996 108684 184664 108712
rect 100996 108672 101002 108684
rect 184658 108672 184664 108684
rect 184716 108672 184722 108724
rect 410794 108672 410800 108724
rect 410852 108712 410858 108724
rect 505922 108712 505928 108724
rect 410852 108684 505928 108712
rect 410852 108672 410858 108684
rect 505922 108672 505928 108684
rect 505980 108672 505986 108724
rect 68370 108604 68376 108656
rect 68428 108644 68434 108656
rect 181898 108644 181904 108656
rect 68428 108616 181904 108644
rect 68428 108604 68434 108616
rect 181898 108604 181904 108616
rect 181956 108604 181962 108656
rect 412542 108604 412548 108656
rect 412600 108644 412606 108656
rect 416130 108644 416136 108656
rect 412600 108616 416136 108644
rect 412600 108604 412606 108616
rect 416130 108604 416136 108616
rect 416188 108604 416194 108656
rect 418890 108604 418896 108656
rect 418948 108644 418954 108656
rect 520918 108644 520924 108656
rect 418948 108616 520924 108644
rect 418948 108604 418954 108616
rect 520918 108604 520924 108616
rect 520976 108604 520982 108656
rect 61102 108536 61108 108588
rect 61160 108576 61166 108588
rect 181714 108576 181720 108588
rect 61160 108548 181720 108576
rect 61160 108536 61166 108548
rect 181714 108536 181720 108548
rect 181772 108536 181778 108588
rect 410886 108536 410892 108588
rect 410944 108576 410950 108588
rect 513374 108576 513380 108588
rect 410944 108548 513380 108576
rect 410944 108536 410950 108548
rect 513374 108536 513380 108548
rect 513432 108536 513438 108588
rect 56042 108468 56048 108520
rect 56100 108508 56106 108520
rect 181990 108508 181996 108520
rect 56100 108480 181996 108508
rect 56100 108468 56106 108480
rect 181990 108468 181996 108480
rect 182048 108468 182054 108520
rect 410978 108468 410984 108520
rect 411036 108508 411042 108520
rect 515858 108508 515864 108520
rect 411036 108480 515864 108508
rect 411036 108468 411042 108480
rect 515858 108468 515864 108480
rect 515916 108468 515922 108520
rect 53650 108400 53656 108452
rect 53708 108440 53714 108452
rect 184106 108440 184112 108452
rect 53708 108412 184112 108440
rect 53708 108400 53714 108412
rect 184106 108400 184112 108412
rect 184164 108400 184170 108452
rect 411070 108400 411076 108452
rect 411128 108440 411134 108452
rect 518434 108440 518440 108452
rect 411128 108412 518440 108440
rect 411128 108400 411134 108412
rect 518434 108400 518440 108412
rect 518492 108400 518498 108452
rect 50798 108332 50804 108384
rect 50856 108372 50862 108384
rect 184566 108372 184572 108384
rect 50856 108344 184572 108372
rect 50856 108332 50862 108344
rect 184566 108332 184572 108344
rect 184624 108332 184630 108384
rect 413278 108332 413284 108384
rect 413336 108372 413342 108384
rect 525886 108372 525892 108384
rect 413336 108344 525892 108372
rect 413336 108332 413342 108344
rect 525886 108332 525892 108344
rect 525944 108332 525950 108384
rect 48314 108264 48320 108316
rect 48372 108304 48378 108316
rect 187234 108304 187240 108316
rect 48372 108276 187240 108304
rect 48372 108264 48378 108276
rect 187234 108264 187240 108276
rect 187292 108264 187298 108316
rect 285674 108264 285680 108316
rect 285732 108304 285738 108316
rect 358814 108304 358820 108316
rect 285732 108276 358820 108304
rect 285732 108264 285738 108276
rect 358814 108264 358820 108276
rect 358872 108264 358878 108316
rect 388622 108264 388628 108316
rect 388680 108304 388686 108316
rect 523310 108304 523316 108316
rect 388680 108276 523316 108304
rect 388680 108264 388686 108276
rect 523310 108264 523316 108276
rect 523368 108264 523374 108316
rect 414382 108196 414388 108248
rect 414440 108236 414446 108248
rect 414842 108236 414848 108248
rect 414440 108208 414848 108236
rect 414440 108196 414446 108208
rect 414842 108196 414848 108208
rect 414900 108236 414906 108248
rect 414900 108208 422294 108236
rect 414900 108196 414906 108208
rect 415118 108128 415124 108180
rect 415176 108168 415182 108180
rect 416406 108168 416412 108180
rect 415176 108140 416412 108168
rect 415176 108128 415182 108140
rect 416406 108128 416412 108140
rect 416464 108128 416470 108180
rect 18414 108060 18420 108112
rect 18472 108100 18478 108112
rect 19242 108100 19248 108112
rect 18472 108072 19248 108100
rect 18472 108060 18478 108072
rect 19242 108060 19248 108072
rect 19300 108060 19306 108112
rect 19518 107992 19524 108044
rect 19576 108032 19582 108044
rect 19794 108032 19800 108044
rect 19576 108004 19800 108032
rect 19576 107992 19582 108004
rect 19794 107992 19800 108004
rect 19852 107992 19858 108044
rect 414566 107992 414572 108044
rect 414624 108032 414630 108044
rect 415210 108032 415216 108044
rect 414624 108004 415216 108032
rect 414624 107992 414630 108004
rect 415210 107992 415216 108004
rect 415268 107992 415274 108044
rect 422266 108032 422294 108208
rect 457990 108032 457996 108044
rect 422266 108004 457996 108032
rect 457990 107992 457996 108004
rect 458048 107992 458054 108044
rect 418062 107924 418068 107976
rect 418120 107964 418126 107976
rect 418430 107964 418436 107976
rect 418120 107936 418436 107964
rect 418120 107924 418126 107936
rect 418430 107924 418436 107936
rect 418488 107964 418494 107976
rect 452562 107964 452568 107976
rect 418488 107936 452568 107964
rect 418488 107924 418494 107936
rect 452562 107924 452568 107936
rect 452620 107924 452626 107976
rect 418338 107856 418344 107908
rect 418396 107896 418402 107908
rect 419258 107896 419264 107908
rect 418396 107868 419264 107896
rect 418396 107856 418402 107868
rect 419258 107856 419264 107868
rect 419316 107896 419322 107908
rect 456978 107896 456984 107908
rect 419316 107868 456984 107896
rect 419316 107856 419322 107868
rect 456978 107856 456984 107868
rect 457036 107856 457042 107908
rect 19242 107788 19248 107840
rect 19300 107828 19306 107840
rect 19300 107800 26234 107828
rect 19300 107788 19306 107800
rect 16482 107720 16488 107772
rect 16540 107760 16546 107772
rect 19610 107760 19616 107772
rect 16540 107732 19616 107760
rect 16540 107720 16546 107732
rect 19610 107720 19616 107732
rect 19668 107760 19674 107772
rect 19668 107732 20668 107760
rect 19668 107720 19674 107732
rect 18690 107584 18696 107636
rect 18748 107624 18754 107636
rect 19426 107624 19432 107636
rect 18748 107596 19432 107624
rect 18748 107584 18754 107596
rect 19426 107584 19432 107596
rect 19484 107584 19490 107636
rect 20640 107624 20668 107732
rect 26206 107692 26234 107800
rect 416406 107788 416412 107840
rect 416464 107828 416470 107840
rect 455782 107828 455788 107840
rect 416464 107800 455788 107828
rect 416464 107788 416470 107800
rect 455782 107788 455788 107800
rect 455840 107788 455846 107840
rect 416130 107720 416136 107772
rect 416188 107760 416194 107772
rect 458174 107760 458180 107772
rect 416188 107732 458180 107760
rect 416188 107720 416194 107732
rect 458174 107720 458180 107732
rect 458232 107720 458238 107772
rect 50154 107692 50160 107704
rect 26206 107664 50160 107692
rect 50154 107652 50160 107664
rect 50212 107652 50218 107704
rect 416314 107652 416320 107704
rect 416372 107692 416378 107704
rect 418154 107692 418160 107704
rect 416372 107664 418160 107692
rect 416372 107652 416378 107664
rect 418154 107652 418160 107664
rect 418212 107692 418218 107704
rect 418890 107692 418896 107704
rect 418212 107664 418896 107692
rect 418212 107652 418218 107664
rect 418890 107652 418896 107664
rect 418948 107652 418954 107704
rect 456978 107652 456984 107704
rect 457036 107692 457042 107704
rect 457036 107664 471928 107692
rect 457036 107652 457042 107664
rect 59630 107624 59636 107636
rect 20640 107596 59636 107624
rect 59630 107584 59636 107596
rect 59688 107584 59694 107636
rect 63586 107584 63592 107636
rect 63644 107624 63650 107636
rect 191190 107624 191196 107636
rect 63644 107596 191196 107624
rect 63644 107584 63650 107596
rect 191190 107584 191196 107596
rect 191248 107584 191254 107636
rect 392578 107584 392584 107636
rect 392636 107624 392642 107636
rect 450630 107624 450636 107636
rect 392636 107596 450636 107624
rect 392636 107584 392642 107596
rect 450630 107584 450636 107596
rect 450688 107584 450694 107636
rect 458174 107584 458180 107636
rect 458232 107624 458238 107636
rect 459462 107624 459468 107636
rect 458232 107596 459468 107624
rect 458232 107584 458238 107596
rect 459462 107584 459468 107596
rect 459520 107624 459526 107636
rect 471900 107624 471928 107664
rect 475654 107624 475660 107636
rect 459520 107596 470594 107624
rect 471900 107596 475660 107624
rect 459520 107584 459526 107596
rect 19058 107516 19064 107568
rect 19116 107556 19122 107568
rect 36906 107556 36912 107568
rect 19116 107528 36912 107556
rect 19116 107516 19122 107528
rect 36906 107516 36912 107528
rect 36964 107516 36970 107568
rect 50154 107516 50160 107568
rect 50212 107556 50218 107568
rect 68646 107556 68652 107568
rect 50212 107528 68652 107556
rect 50212 107516 50218 107528
rect 68646 107516 68652 107528
rect 68704 107516 68710 107568
rect 73706 107516 73712 107568
rect 73764 107556 73770 107568
rect 186958 107556 186964 107568
rect 73764 107528 186964 107556
rect 73764 107516 73770 107528
rect 186958 107516 186964 107528
rect 187016 107516 187022 107568
rect 408126 107516 408132 107568
rect 408184 107556 408190 107568
rect 458358 107556 458364 107568
rect 408184 107528 458364 107556
rect 408184 107516 408190 107528
rect 458358 107516 458364 107528
rect 458416 107516 458422 107568
rect 470566 107556 470594 107596
rect 475654 107584 475660 107596
rect 475712 107584 475718 107636
rect 478046 107556 478052 107568
rect 470566 107528 478052 107556
rect 478046 107516 478052 107528
rect 478104 107516 478110 107568
rect 18506 107448 18512 107500
rect 18564 107488 18570 107500
rect 19610 107488 19616 107500
rect 18564 107460 19616 107488
rect 18564 107448 18570 107460
rect 19610 107448 19616 107460
rect 19668 107448 19674 107500
rect 43162 107488 43168 107500
rect 41524 107460 43168 107488
rect 16114 107380 16120 107432
rect 16172 107420 16178 107432
rect 18782 107420 18788 107432
rect 16172 107392 18788 107420
rect 16172 107380 16178 107392
rect 18782 107380 18788 107392
rect 18840 107380 18846 107432
rect 18966 107380 18972 107432
rect 19024 107420 19030 107432
rect 35894 107420 35900 107432
rect 19024 107392 35900 107420
rect 19024 107380 19030 107392
rect 35894 107380 35900 107392
rect 35952 107380 35958 107432
rect 19150 107312 19156 107364
rect 19208 107352 19214 107364
rect 38102 107352 38108 107364
rect 19208 107324 38108 107352
rect 19208 107312 19214 107324
rect 38102 107312 38108 107324
rect 38160 107312 38166 107364
rect 18874 107244 18880 107296
rect 18932 107284 18938 107296
rect 39574 107284 39580 107296
rect 18932 107256 39580 107284
rect 18932 107244 18938 107256
rect 39574 107244 39580 107256
rect 39632 107244 39638 107296
rect 19702 107176 19708 107228
rect 19760 107216 19766 107228
rect 41524 107216 41552 107460
rect 43162 107448 43168 107460
rect 43220 107488 43226 107500
rect 61654 107488 61660 107500
rect 43220 107460 61660 107488
rect 43220 107448 43226 107460
rect 61654 107448 61660 107460
rect 61712 107448 61718 107500
rect 61746 107448 61752 107500
rect 61804 107488 61810 107500
rect 75638 107488 75644 107500
rect 61804 107460 75644 107488
rect 61804 107448 61810 107460
rect 75638 107448 75644 107460
rect 75696 107448 75702 107500
rect 76098 107448 76104 107500
rect 76156 107488 76162 107500
rect 187142 107488 187148 107500
rect 76156 107460 187148 107488
rect 76156 107448 76162 107460
rect 187142 107448 187148 107460
rect 187200 107448 187206 107500
rect 408034 107448 408040 107500
rect 408092 107488 408098 107500
rect 455966 107488 455972 107500
rect 408092 107460 455972 107488
rect 408092 107448 408098 107460
rect 455966 107448 455972 107460
rect 456024 107448 456030 107500
rect 474366 107488 474372 107500
rect 456076 107460 474372 107488
rect 52270 107380 52276 107432
rect 52328 107420 52334 107432
rect 69750 107420 69756 107432
rect 52328 107392 69756 107420
rect 52328 107380 52334 107392
rect 69750 107380 69756 107392
rect 69808 107380 69814 107432
rect 78490 107380 78496 107432
rect 78548 107420 78554 107432
rect 187050 107420 187056 107432
rect 78548 107392 187056 107420
rect 78548 107380 78554 107392
rect 187050 107380 187056 107392
rect 187108 107380 187114 107432
rect 417878 107380 417884 107432
rect 417936 107420 417942 107432
rect 419258 107420 419264 107432
rect 417936 107392 419264 107420
rect 417936 107380 417942 107392
rect 419258 107380 419264 107392
rect 419316 107380 419322 107432
rect 455782 107380 455788 107432
rect 455840 107420 455846 107432
rect 456076 107420 456104 107460
rect 474366 107448 474372 107460
rect 474424 107448 474430 107500
rect 471146 107420 471152 107432
rect 455840 107392 456104 107420
rect 460906 107392 471152 107420
rect 455840 107380 455846 107392
rect 44358 107312 44364 107364
rect 44416 107352 44422 107364
rect 45370 107352 45376 107364
rect 44416 107324 45376 107352
rect 44416 107312 44422 107324
rect 45370 107312 45376 107324
rect 45428 107352 45434 107364
rect 63862 107352 63868 107364
rect 45428 107324 63868 107352
rect 45428 107312 45434 107324
rect 63862 107312 63868 107324
rect 63920 107312 63926 107364
rect 86034 107312 86040 107364
rect 86092 107352 86098 107364
rect 158162 107352 158168 107364
rect 86092 107324 158168 107352
rect 86092 107312 86098 107324
rect 158162 107312 158168 107324
rect 158220 107312 158226 107364
rect 418890 107312 418896 107364
rect 418948 107352 418954 107364
rect 418948 107324 451274 107352
rect 418948 107312 418954 107324
rect 46566 107244 46572 107296
rect 46624 107284 46630 107296
rect 65150 107284 65156 107296
rect 46624 107256 65156 107284
rect 46624 107244 46630 107256
rect 65150 107244 65156 107256
rect 65208 107244 65214 107296
rect 88242 107244 88248 107296
rect 88300 107284 88306 107296
rect 156598 107284 156604 107296
rect 88300 107256 156604 107284
rect 88300 107244 88306 107256
rect 156598 107244 156604 107256
rect 156656 107244 156662 107296
rect 44266 107216 44272 107228
rect 19760 107188 41552 107216
rect 44100 107188 44272 107216
rect 19760 107176 19766 107188
rect 19518 107108 19524 107160
rect 19576 107148 19582 107160
rect 44100 107148 44128 107188
rect 44266 107176 44272 107188
rect 44324 107176 44330 107228
rect 48774 107176 48780 107228
rect 48832 107216 48838 107228
rect 67634 107216 67640 107228
rect 48832 107188 67640 107216
rect 48832 107176 48838 107188
rect 67634 107176 67640 107188
rect 67692 107176 67698 107228
rect 93578 107176 93584 107228
rect 93636 107216 93642 107228
rect 158070 107216 158076 107228
rect 93636 107188 158076 107216
rect 93636 107176 93642 107188
rect 158070 107176 158076 107188
rect 158128 107176 158134 107228
rect 418706 107176 418712 107228
rect 418764 107216 418770 107228
rect 436094 107216 436100 107228
rect 418764 107188 436100 107216
rect 418764 107176 418770 107188
rect 436094 107176 436100 107188
rect 436152 107176 436158 107228
rect 451246 107216 451274 107324
rect 452562 107312 452568 107364
rect 452620 107352 452626 107364
rect 460906 107352 460934 107392
rect 471146 107380 471152 107392
rect 471204 107380 471210 107432
rect 452620 107324 460934 107352
rect 452620 107312 452626 107324
rect 452470 107244 452476 107296
rect 452528 107284 452534 107296
rect 469766 107284 469772 107296
rect 452528 107256 469772 107284
rect 452528 107244 452534 107256
rect 469766 107244 469772 107256
rect 469824 107244 469830 107296
rect 459554 107216 459560 107228
rect 451246 107188 459560 107216
rect 459554 107176 459560 107188
rect 459612 107176 459618 107228
rect 19576 107120 44128 107148
rect 19576 107108 19582 107120
rect 44174 107108 44180 107160
rect 44232 107148 44238 107160
rect 47578 107148 47584 107160
rect 44232 107120 47584 107148
rect 44232 107108 44238 107120
rect 47578 107108 47584 107120
rect 47636 107148 47642 107160
rect 66254 107148 66260 107160
rect 47636 107120 66260 107148
rect 47636 107108 47642 107120
rect 66254 107108 66260 107120
rect 66312 107108 66318 107160
rect 120994 107108 121000 107160
rect 121052 107148 121058 107160
rect 181806 107148 181812 107160
rect 121052 107120 181812 107148
rect 121052 107108 121058 107120
rect 181806 107108 181812 107120
rect 181864 107108 181870 107160
rect 419810 107108 419816 107160
rect 419868 107148 419874 107160
rect 438118 107148 438124 107160
rect 419868 107120 438124 107148
rect 419868 107108 419874 107120
rect 438118 107108 438124 107120
rect 438176 107108 438182 107160
rect 444282 107108 444288 107160
rect 444340 107148 444346 107160
rect 461670 107148 461676 107160
rect 444340 107120 461676 107148
rect 444340 107108 444346 107120
rect 461670 107108 461676 107120
rect 461728 107108 461734 107160
rect 17126 107040 17132 107092
rect 17184 107080 17190 107092
rect 52362 107080 52368 107092
rect 17184 107052 52368 107080
rect 17184 107040 17190 107052
rect 52362 107040 52368 107052
rect 52420 107080 52426 107092
rect 52420 107052 54708 107080
rect 52420 107040 52426 107052
rect 15562 106972 15568 107024
rect 15620 107012 15626 107024
rect 16206 107012 16212 107024
rect 15620 106984 16212 107012
rect 15620 106972 15626 106984
rect 16206 106972 16212 106984
rect 16264 107012 16270 107024
rect 51258 107012 51264 107024
rect 16264 106984 51264 107012
rect 16264 106972 16270 106984
rect 51258 106972 51264 106984
rect 51316 107012 51322 107024
rect 52270 107012 52276 107024
rect 51316 106984 52276 107012
rect 51316 106972 51322 106984
rect 52270 106972 52276 106984
rect 52328 106972 52334 107024
rect 54680 107012 54708 107052
rect 59354 107040 59360 107092
rect 59412 107080 59418 107092
rect 60550 107080 60556 107092
rect 59412 107052 60556 107080
rect 59412 107040 59418 107052
rect 60550 107040 60556 107052
rect 60608 107080 60614 107092
rect 79134 107080 79140 107092
rect 60608 107052 79140 107080
rect 60608 107040 60614 107052
rect 79134 107040 79140 107052
rect 79192 107040 79198 107092
rect 123386 107040 123392 107092
rect 123444 107080 123450 107092
rect 181622 107080 181628 107092
rect 123444 107052 181628 107080
rect 123444 107040 123450 107052
rect 181622 107040 181628 107052
rect 181680 107040 181686 107092
rect 419718 107040 419724 107092
rect 419776 107080 419782 107092
rect 439590 107080 439596 107092
rect 419776 107052 439596 107080
rect 419776 107040 419782 107052
rect 439590 107040 439596 107052
rect 439648 107040 439654 107092
rect 444190 107080 444196 107092
rect 441586 107052 444196 107080
rect 71222 107012 71228 107024
rect 54680 106984 71228 107012
rect 71222 106972 71228 106984
rect 71280 106972 71286 107024
rect 98546 106972 98552 107024
rect 98604 107012 98610 107024
rect 156690 107012 156696 107024
rect 98604 106984 156696 107012
rect 98604 106972 98610 106984
rect 156690 106972 156696 106984
rect 156748 106972 156754 107024
rect 339494 106972 339500 107024
rect 339552 107012 339558 107024
rect 359642 107012 359648 107024
rect 339552 106984 359648 107012
rect 339552 106972 339558 106984
rect 359642 106972 359648 106984
rect 359700 106972 359706 107024
rect 415118 106972 415124 107024
rect 415176 107012 415182 107024
rect 441586 107012 441614 107052
rect 444190 107040 444196 107052
rect 444248 107080 444254 107092
rect 462774 107080 462780 107092
rect 444248 107052 462780 107080
rect 444248 107040 444254 107052
rect 462774 107040 462780 107052
rect 462832 107040 462838 107092
rect 454586 107012 454592 107024
rect 415176 106984 441614 107012
rect 451246 106984 454592 107012
rect 415176 106972 415182 106984
rect 15010 106904 15016 106956
rect 15068 106944 15074 106956
rect 53466 106944 53472 106956
rect 15068 106916 53472 106944
rect 15068 106904 15074 106916
rect 53466 106904 53472 106916
rect 53524 106944 53530 106956
rect 72142 106944 72148 106956
rect 53524 106916 72148 106944
rect 53524 106904 53530 106916
rect 72142 106904 72148 106916
rect 72200 106904 72206 106956
rect 335354 106904 335360 106956
rect 335412 106944 335418 106956
rect 418890 106944 418896 106956
rect 335412 106916 418896 106944
rect 335412 106904 335418 106916
rect 418890 106904 418896 106916
rect 418948 106904 418954 106956
rect 419902 106904 419908 106956
rect 419960 106944 419966 106956
rect 451246 106944 451274 106984
rect 454586 106972 454592 106984
rect 454644 107012 454650 107024
rect 473354 107012 473360 107024
rect 454644 106984 473360 107012
rect 454644 106972 454650 106984
rect 473354 106972 473360 106984
rect 473412 106972 473418 107024
rect 419960 106916 451274 106944
rect 419960 106904 419966 106916
rect 459554 106904 459560 106956
rect 459612 106944 459618 106956
rect 460658 106944 460664 106956
rect 459612 106916 460664 106944
rect 459612 106904 459618 106916
rect 460658 106904 460664 106916
rect 460716 106944 460722 106956
rect 479150 106944 479156 106956
rect 460716 106916 479156 106944
rect 460716 106904 460722 106916
rect 479150 106904 479156 106916
rect 479208 106904 479214 106956
rect 59630 106836 59636 106888
rect 59688 106876 59694 106888
rect 77662 106876 77668 106888
rect 59688 106848 77668 106876
rect 59688 106836 59694 106848
rect 77662 106836 77668 106848
rect 77720 106836 77726 106888
rect 418982 106836 418988 106888
rect 419040 106876 419046 106888
rect 419350 106876 419356 106888
rect 419040 106848 419356 106876
rect 419040 106836 419046 106848
rect 419350 106836 419356 106848
rect 419408 106876 419414 106888
rect 437014 106876 437020 106888
rect 419408 106848 437020 106876
rect 419408 106836 419414 106848
rect 437014 106836 437020 106848
rect 437072 106836 437078 106888
rect 44266 106768 44272 106820
rect 44324 106808 44330 106820
rect 62574 106808 62580 106820
rect 44324 106780 62580 106808
rect 44324 106768 44330 106780
rect 62574 106768 62580 106780
rect 62632 106768 62638 106820
rect 410610 106768 410616 106820
rect 410668 106808 410674 106820
rect 453574 106808 453580 106820
rect 410668 106780 453580 106808
rect 410668 106768 410674 106780
rect 453574 106768 453580 106780
rect 453632 106768 453638 106820
rect 448514 106632 448520 106684
rect 448572 106672 448578 106684
rect 467006 106672 467012 106684
rect 448572 106644 467012 106672
rect 448572 106632 448578 106644
rect 467006 106632 467012 106644
rect 467064 106632 467070 106684
rect 447134 106564 447140 106616
rect 447192 106604 447198 106616
rect 465718 106604 465724 106616
rect 447192 106576 465724 106604
rect 447192 106564 447198 106576
rect 465718 106564 465724 106576
rect 465776 106564 465782 106616
rect 19794 106496 19800 106548
rect 19852 106536 19858 106548
rect 40494 106536 40500 106548
rect 19852 106508 40500 106536
rect 19852 106496 19858 106508
rect 40494 106496 40500 106508
rect 40552 106496 40558 106548
rect 42794 106496 42800 106548
rect 42852 106536 42858 106548
rect 48774 106536 48780 106548
rect 42852 106508 48780 106536
rect 42852 106496 42858 106508
rect 48774 106496 48780 106508
rect 48832 106496 48838 106548
rect 449894 106496 449900 106548
rect 449952 106536 449958 106548
rect 468662 106536 468668 106548
rect 449952 106508 468668 106536
rect 449952 106496 449958 106508
rect 468662 106496 468668 106508
rect 468720 106496 468726 106548
rect 18322 106428 18328 106480
rect 18380 106468 18386 106480
rect 18782 106468 18788 106480
rect 18380 106440 18788 106468
rect 18380 106428 18386 106440
rect 18782 106428 18788 106440
rect 18840 106468 18846 106480
rect 44358 106468 44364 106480
rect 18840 106440 44364 106468
rect 18840 106428 18846 106440
rect 44358 106428 44364 106440
rect 44416 106428 44422 106480
rect 55766 106428 55772 106480
rect 55824 106468 55830 106480
rect 74350 106468 74356 106480
rect 55824 106440 74356 106468
rect 55824 106428 55830 106440
rect 74350 106428 74356 106440
rect 74408 106428 74414 106480
rect 418062 106428 418068 106480
rect 418120 106468 418126 106480
rect 440510 106468 440516 106480
rect 418120 106440 440516 106468
rect 418120 106428 418126 106440
rect 440510 106428 440516 106440
rect 440568 106428 440574 106480
rect 445662 106428 445668 106480
rect 445720 106468 445726 106480
rect 463878 106468 463884 106480
rect 445720 106440 463884 106468
rect 445720 106428 445726 106440
rect 463878 106428 463884 106440
rect 463936 106428 463942 106480
rect 19426 106360 19432 106412
rect 19484 106400 19490 106412
rect 46566 106400 46572 106412
rect 19484 106372 46572 106400
rect 19484 106360 19490 106372
rect 46566 106360 46572 106372
rect 46624 106360 46630 106412
rect 55306 106360 55312 106412
rect 55364 106400 55370 106412
rect 73246 106400 73252 106412
rect 55364 106372 73252 106400
rect 55364 106360 55370 106372
rect 73246 106360 73252 106372
rect 73304 106360 73310 106412
rect 417050 106360 417056 106412
rect 417108 106400 417114 106412
rect 441614 106400 441620 106412
rect 417108 106372 441620 106400
rect 417108 106360 417114 106372
rect 441614 106360 441620 106372
rect 441672 106360 441678 106412
rect 446398 106360 446404 106412
rect 446456 106400 446462 106412
rect 465166 106400 465172 106412
rect 446456 106372 465172 106400
rect 446456 106360 446462 106372
rect 465166 106360 465172 106372
rect 465224 106360 465230 106412
rect 19610 106292 19616 106344
rect 19668 106332 19674 106344
rect 59354 106332 59360 106344
rect 19668 106304 59360 106332
rect 19668 106292 19674 106304
rect 59354 106292 59360 106304
rect 59412 106292 59418 106344
rect 419258 106292 419264 106344
rect 419316 106332 419322 106344
rect 443086 106332 443092 106344
rect 419316 106304 443092 106332
rect 419316 106292 419322 106304
rect 443086 106292 443092 106304
rect 443144 106332 443150 106344
rect 444282 106332 444288 106344
rect 443144 106304 444288 106332
rect 443144 106292 443150 106304
rect 444282 106292 444288 106304
rect 444340 106292 444346 106344
rect 453942 106292 453948 106344
rect 454000 106332 454006 106344
rect 472066 106332 472072 106344
rect 454000 106304 472072 106332
rect 454000 106292 454006 106304
rect 472066 106292 472072 106304
rect 472124 106292 472130 106344
rect 17218 106224 17224 106276
rect 17276 106264 17282 106276
rect 150802 106264 150808 106276
rect 17276 106236 150808 106264
rect 17276 106224 17282 106236
rect 150802 106224 150808 106236
rect 150860 106264 150866 106276
rect 157334 106264 157340 106276
rect 150860 106236 157340 106264
rect 150860 106224 150866 106236
rect 157334 106224 157340 106236
rect 157392 106264 157398 106276
rect 351178 106264 351184 106276
rect 157392 106236 351184 106264
rect 157392 106224 157398 106236
rect 351178 106224 351184 106236
rect 351236 106224 351242 106276
rect 415026 106224 415032 106276
rect 415084 106264 415090 106276
rect 416222 106264 416228 106276
rect 415084 106236 416228 106264
rect 415084 106224 415090 106236
rect 416222 106224 416228 106236
rect 416280 106224 416286 106276
rect 417786 106224 417792 106276
rect 417844 106264 417850 106276
rect 550726 106264 550732 106276
rect 417844 106236 550732 106264
rect 417844 106224 417850 106236
rect 550726 106224 550732 106236
rect 550784 106264 550790 106276
rect 557534 106264 557540 106276
rect 550784 106236 557540 106264
rect 550784 106224 550790 106236
rect 557534 106224 557540 106236
rect 557592 106224 557598 106276
rect 14826 106156 14832 106208
rect 14884 106196 14890 106208
rect 15102 106196 15108 106208
rect 14884 106168 15108 106196
rect 14884 106156 14890 106168
rect 15102 106156 15108 106168
rect 15160 106196 15166 106208
rect 44174 106196 44180 106208
rect 15160 106168 44180 106196
rect 15160 106156 15166 106168
rect 44174 106156 44180 106168
rect 44232 106156 44238 106208
rect 414474 106156 414480 106208
rect 414532 106196 414538 106208
rect 415302 106196 415308 106208
rect 414532 106168 415308 106196
rect 414532 106156 414538 106168
rect 415302 106156 415308 106168
rect 415360 106156 415366 106208
rect 417694 106156 417700 106208
rect 417752 106196 417758 106208
rect 418614 106196 418620 106208
rect 417752 106168 418620 106196
rect 417752 106156 417758 106168
rect 418614 106156 418620 106168
rect 418672 106156 418678 106208
rect 419994 106156 420000 106208
rect 420052 106196 420058 106208
rect 453942 106196 453948 106208
rect 420052 106168 453948 106196
rect 420052 106156 420058 106168
rect 453942 106156 453948 106168
rect 454000 106156 454006 106208
rect 16022 106088 16028 106140
rect 16080 106128 16086 106140
rect 16390 106128 16396 106140
rect 16080 106100 16396 106128
rect 16080 106088 16086 106100
rect 16390 106088 16396 106100
rect 16448 106128 16454 106140
rect 42794 106128 42800 106140
rect 16448 106100 42800 106128
rect 16448 106088 16454 106100
rect 42794 106088 42800 106100
rect 42852 106088 42858 106140
rect 415320 106128 415348 106156
rect 447134 106128 447140 106140
rect 415320 106100 447140 106128
rect 447134 106088 447140 106100
rect 447192 106088 447198 106140
rect 414750 106020 414756 106072
rect 414808 106060 414814 106072
rect 446398 106060 446404 106072
rect 414808 106032 446404 106060
rect 414808 106020 414814 106032
rect 446398 106020 446404 106032
rect 446456 106020 446462 106072
rect 219158 105952 219164 106004
rect 219216 105992 219222 106004
rect 251174 105992 251180 106004
rect 219216 105964 251180 105992
rect 219216 105952 219222 105964
rect 251174 105952 251180 105964
rect 251232 105952 251238 106004
rect 280154 105952 280160 106004
rect 280212 105992 280218 106004
rect 357250 105992 357256 106004
rect 280212 105964 357256 105992
rect 280212 105952 280218 105964
rect 357250 105952 357256 105964
rect 357308 105952 357314 106004
rect 414566 105952 414572 106004
rect 414624 105992 414630 106004
rect 445662 105992 445668 106004
rect 414624 105964 445668 105992
rect 414624 105952 414630 105964
rect 445662 105952 445668 105964
rect 445720 105952 445726 106004
rect 219986 105884 219992 105936
rect 220044 105924 220050 105936
rect 252554 105924 252560 105936
rect 220044 105896 252560 105924
rect 220044 105884 220050 105896
rect 252554 105884 252560 105896
rect 252612 105884 252618 105936
rect 278774 105884 278780 105936
rect 278832 105924 278838 105936
rect 357894 105924 357900 105936
rect 278832 105896 357900 105924
rect 278832 105884 278838 105896
rect 357894 105884 357900 105896
rect 357952 105884 357958 105936
rect 219250 105816 219256 105868
rect 219308 105856 219314 105868
rect 255314 105856 255320 105868
rect 219308 105828 255320 105856
rect 219308 105816 219314 105828
rect 255314 105816 255320 105828
rect 255372 105816 255378 105868
rect 277394 105816 277400 105868
rect 277452 105856 277458 105868
rect 357710 105856 357716 105868
rect 277452 105828 357716 105856
rect 277452 105816 277458 105828
rect 357710 105816 357716 105828
rect 357768 105816 357774 105868
rect 217226 105748 217232 105800
rect 217284 105788 217290 105800
rect 259454 105788 259460 105800
rect 217284 105760 259460 105788
rect 217284 105748 217290 105760
rect 259454 105748 259460 105760
rect 259512 105748 259518 105800
rect 274634 105748 274640 105800
rect 274692 105788 274698 105800
rect 357802 105788 357808 105800
rect 274692 105760 357808 105788
rect 274692 105748 274698 105760
rect 357802 105748 357808 105760
rect 357860 105748 357866 105800
rect 15654 105680 15660 105732
rect 15712 105720 15718 105732
rect 18598 105720 18604 105732
rect 15712 105692 18604 105720
rect 15712 105680 15718 105692
rect 18598 105680 18604 105692
rect 18656 105720 18662 105732
rect 55306 105720 55312 105732
rect 18656 105692 55312 105720
rect 18656 105680 18662 105692
rect 55306 105680 55312 105692
rect 55364 105680 55370 105732
rect 216214 105680 216220 105732
rect 216272 105720 216278 105732
rect 262214 105720 262220 105732
rect 216272 105692 262220 105720
rect 216272 105680 216278 105692
rect 262214 105680 262220 105692
rect 262272 105680 262278 105732
rect 273254 105680 273260 105732
rect 273312 105720 273318 105732
rect 357066 105720 357072 105732
rect 273312 105692 357072 105720
rect 273312 105680 273318 105692
rect 357066 105680 357072 105692
rect 357124 105680 357130 105732
rect 15838 105612 15844 105664
rect 15896 105652 15902 105664
rect 18506 105652 18512 105664
rect 15896 105624 18512 105652
rect 15896 105612 15902 105624
rect 18506 105612 18512 105624
rect 18564 105652 18570 105664
rect 55766 105652 55772 105664
rect 18564 105624 55772 105652
rect 18564 105612 18570 105624
rect 55766 105612 55772 105624
rect 55824 105612 55830 105664
rect 216306 105612 216312 105664
rect 216364 105652 216370 105664
rect 263594 105652 263600 105664
rect 216364 105624 263600 105652
rect 216364 105612 216370 105624
rect 263594 105612 263600 105624
rect 263652 105612 263658 105664
rect 270494 105612 270500 105664
rect 270552 105652 270558 105664
rect 358906 105652 358912 105664
rect 270552 105624 358912 105652
rect 270552 105612 270558 105624
rect 358906 105612 358912 105624
rect 358964 105612 358970 105664
rect 418614 105612 418620 105664
rect 418672 105652 418678 105664
rect 449894 105652 449900 105664
rect 418672 105624 449900 105652
rect 418672 105612 418678 105624
rect 449894 105612 449900 105624
rect 449952 105612 449958 105664
rect 16298 105544 16304 105596
rect 16356 105584 16362 105596
rect 18690 105584 18696 105596
rect 16356 105556 18696 105584
rect 16356 105544 16362 105556
rect 18690 105544 18696 105556
rect 18748 105584 18754 105596
rect 57054 105584 57060 105596
rect 18748 105556 57060 105584
rect 18748 105544 18754 105556
rect 57054 105544 57060 105556
rect 57112 105544 57118 105596
rect 218974 105544 218980 105596
rect 219032 105584 219038 105596
rect 266354 105584 266360 105596
rect 219032 105556 266360 105584
rect 219032 105544 219038 105556
rect 266354 105544 266360 105556
rect 266412 105544 266418 105596
rect 269114 105544 269120 105596
rect 269172 105584 269178 105596
rect 358998 105584 359004 105596
rect 269172 105556 359004 105584
rect 269172 105544 269178 105556
rect 358998 105544 359004 105556
rect 359056 105544 359062 105596
rect 414382 105544 414388 105596
rect 414440 105584 414446 105596
rect 414750 105584 414756 105596
rect 414440 105556 414756 105584
rect 414440 105544 414446 105556
rect 414750 105544 414756 105556
rect 414808 105544 414814 105596
rect 416222 105544 416228 105596
rect 416280 105584 416286 105596
rect 448514 105584 448520 105596
rect 416280 105556 448520 105584
rect 416280 105544 416286 105556
rect 448514 105544 448520 105556
rect 448572 105544 448578 105596
rect 17034 104796 17040 104848
rect 17092 104836 17098 104848
rect 390646 104836 390652 104848
rect 17092 104808 390652 104836
rect 17092 104796 17098 104808
rect 390646 104796 390652 104808
rect 390704 104836 390710 104848
rect 417142 104836 417148 104848
rect 390704 104808 417148 104836
rect 390704 104796 390710 104808
rect 417142 104796 417148 104808
rect 417200 104836 417206 104848
rect 417418 104836 417424 104848
rect 417200 104808 417424 104836
rect 417200 104796 417206 104808
rect 417418 104796 417424 104808
rect 417476 104796 417482 104848
rect 219894 104728 219900 104780
rect 219952 104768 219958 104780
rect 222838 104768 222844 104780
rect 219952 104740 222844 104768
rect 219952 104728 219958 104740
rect 222838 104728 222844 104740
rect 222896 104728 222902 104780
rect 219710 104660 219716 104712
rect 219768 104700 219774 104712
rect 228358 104700 228364 104712
rect 219768 104672 228364 104700
rect 219768 104660 219774 104672
rect 228358 104660 228364 104672
rect 228416 104660 228422 104712
rect 351914 104592 351920 104644
rect 351972 104632 351978 104644
rect 411990 104632 411996 104644
rect 351972 104604 411996 104632
rect 351972 104592 351978 104604
rect 411990 104592 411996 104604
rect 412048 104592 412054 104644
rect 350534 104524 350540 104576
rect 350592 104564 350598 104576
rect 414934 104564 414940 104576
rect 350592 104536 414940 104564
rect 350592 104524 350598 104536
rect 414934 104524 414940 104536
rect 414992 104524 414998 104576
rect 219802 104456 219808 104508
rect 219860 104496 219866 104508
rect 223022 104496 223028 104508
rect 219860 104468 223028 104496
rect 219860 104456 219866 104468
rect 223022 104456 223028 104468
rect 223080 104456 223086 104508
rect 349154 104456 349160 104508
rect 349212 104496 349218 104508
rect 414750 104496 414756 104508
rect 349212 104468 414756 104496
rect 349212 104456 349218 104468
rect 414750 104456 414756 104468
rect 414808 104456 414814 104508
rect 346394 104388 346400 104440
rect 346452 104428 346458 104440
rect 414842 104428 414848 104440
rect 346452 104400 414848 104428
rect 346452 104388 346458 104400
rect 414842 104388 414848 104400
rect 414900 104388 414906 104440
rect 219066 104320 219072 104372
rect 219124 104360 219130 104372
rect 225598 104360 225604 104372
rect 219124 104332 225604 104360
rect 219124 104320 219130 104332
rect 225598 104320 225604 104332
rect 225656 104320 225662 104372
rect 284294 104320 284300 104372
rect 284352 104360 284358 104372
rect 359090 104360 359096 104372
rect 284352 104332 359096 104360
rect 284352 104320 284358 104332
rect 359090 104320 359096 104332
rect 359148 104320 359154 104372
rect 282914 104252 282920 104304
rect 282972 104292 282978 104304
rect 359274 104292 359280 104304
rect 282972 104264 359280 104292
rect 282972 104252 282978 104264
rect 359274 104252 359280 104264
rect 359332 104252 359338 104304
rect 217134 104184 217140 104236
rect 217192 104224 217198 104236
rect 225782 104224 225788 104236
rect 217192 104196 225788 104224
rect 217192 104184 217198 104196
rect 225782 104184 225788 104196
rect 225840 104184 225846 104236
rect 281534 104184 281540 104236
rect 281592 104224 281598 104236
rect 359182 104224 359188 104236
rect 281592 104196 359188 104224
rect 281592 104184 281598 104196
rect 359182 104184 359188 104196
rect 359240 104184 359246 104236
rect 218054 104116 218060 104168
rect 218112 104156 218118 104168
rect 231118 104156 231124 104168
rect 218112 104128 231124 104156
rect 218112 104116 218118 104128
rect 231118 104116 231124 104128
rect 231176 104116 231182 104168
rect 329834 104116 329840 104168
rect 329892 104156 329898 104168
rect 418798 104156 418804 104168
rect 329892 104128 418804 104156
rect 329892 104116 329898 104128
rect 418798 104116 418804 104128
rect 418856 104116 418862 104168
rect 216122 103504 216128 103556
rect 216180 103544 216186 103556
rect 359734 103544 359740 103556
rect 216180 103516 359740 103544
rect 216180 103504 216186 103516
rect 359734 103504 359740 103516
rect 359792 103504 359798 103556
rect 183554 102756 183560 102808
rect 183612 102796 183618 102808
rect 219434 102796 219440 102808
rect 183612 102768 219440 102796
rect 183612 102756 183618 102768
rect 219434 102756 219440 102768
rect 219492 102756 219498 102808
rect 360102 99288 360108 99340
rect 360160 99328 360166 99340
rect 387058 99328 387064 99340
rect 360160 99300 387064 99328
rect 360160 99288 360166 99300
rect 387058 99288 387064 99300
rect 387116 99288 387122 99340
rect 356974 98744 356980 98796
rect 357032 98744 357038 98796
rect 158898 98608 158904 98660
rect 158956 98648 158962 98660
rect 170490 98648 170496 98660
rect 158956 98620 170496 98648
rect 158956 98608 158962 98620
rect 170490 98608 170496 98620
rect 170548 98608 170554 98660
rect 356992 98592 357020 98744
rect 357158 98608 357164 98660
rect 357216 98608 357222 98660
rect 356974 98540 356980 98592
rect 357032 98540 357038 98592
rect 357176 98456 357204 98608
rect 357158 98404 357164 98456
rect 357216 98404 357222 98456
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 14550 71720 14556 71732
rect 3384 71692 14556 71720
rect 3384 71680 3390 71692
rect 14550 71680 14556 71692
rect 14608 71680 14614 71732
rect 3326 59304 3332 59356
rect 3384 59344 3390 59356
rect 14458 59344 14464 59356
rect 3384 59316 14464 59344
rect 3384 59304 3390 59316
rect 14458 59304 14464 59316
rect 14516 59304 14522 59356
rect 170490 57876 170496 57928
rect 170548 57916 170554 57928
rect 216122 57916 216128 57928
rect 170548 57888 216128 57916
rect 170548 57876 170554 57888
rect 216122 57876 216128 57888
rect 216180 57916 216186 57928
rect 216674 57916 216680 57928
rect 216180 57888 216680 57916
rect 216180 57876 216186 57888
rect 216674 57876 216680 57888
rect 216732 57876 216738 57928
rect 191558 56516 191564 56568
rect 191616 56556 191622 56568
rect 216674 56556 216680 56568
rect 191616 56528 216680 56556
rect 191616 56516 191622 56528
rect 216674 56516 216680 56528
rect 216732 56516 216738 56568
rect 189810 53728 189816 53780
rect 189868 53768 189874 53780
rect 216674 53768 216680 53780
rect 189868 53740 216680 53768
rect 189868 53728 189874 53740
rect 216674 53728 216680 53740
rect 216732 53728 216738 53780
rect 189718 53660 189724 53712
rect 189776 53700 189782 53712
rect 216766 53700 216772 53712
rect 189776 53672 216772 53700
rect 189776 53660 189782 53672
rect 216766 53660 216772 53672
rect 216824 53660 216830 53712
rect 189902 52368 189908 52420
rect 189960 52408 189966 52420
rect 216766 52408 216772 52420
rect 189960 52380 216772 52408
rect 189960 52368 189966 52380
rect 216766 52368 216772 52380
rect 216824 52368 216830 52420
rect 189994 51008 190000 51060
rect 190052 51048 190058 51060
rect 216674 51048 216680 51060
rect 190052 51020 216680 51048
rect 190052 51008 190058 51020
rect 216674 51008 216680 51020
rect 216732 51008 216738 51060
rect 190086 48220 190092 48272
rect 190144 48260 190150 48272
rect 216674 48260 216680 48272
rect 190144 48232 216680 48260
rect 190144 48220 190150 48232
rect 216674 48220 216680 48232
rect 216732 48220 216738 48272
rect 558178 46860 558184 46912
rect 558236 46900 558242 46912
rect 580166 46900 580172 46912
rect 558236 46872 580172 46900
rect 558236 46860 558242 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3326 45500 3332 45552
rect 3384 45540 3390 45552
rect 7558 45540 7564 45552
rect 3384 45512 7564 45540
rect 3384 45500 3390 45512
rect 7558 45500 7564 45512
rect 7616 45500 7622 45552
rect 3326 33056 3332 33108
rect 3384 33096 3390 33108
rect 19978 33096 19984 33108
rect 3384 33068 19984 33096
rect 3384 33056 3390 33068
rect 19978 33056 19984 33068
rect 20036 33056 20042 33108
rect 391198 28908 391204 28960
rect 391256 28948 391262 28960
rect 416774 28948 416780 28960
rect 391256 28920 416780 28948
rect 391256 28908 391262 28920
rect 416774 28908 416780 28920
rect 416832 28908 416838 28960
rect 371142 28228 371148 28280
rect 371200 28268 371206 28280
rect 416866 28268 416872 28280
rect 371200 28240 416872 28268
rect 371200 28228 371206 28240
rect 416866 28228 416872 28240
rect 416924 28228 416930 28280
rect 418706 22584 418712 22636
rect 418764 22624 418770 22636
rect 419166 22624 419172 22636
rect 418764 22596 419172 22624
rect 418764 22584 418770 22596
rect 419166 22584 419172 22596
rect 419224 22584 419230 22636
rect 418430 22380 418436 22432
rect 418488 22420 418494 22432
rect 418614 22420 418620 22432
rect 418488 22392 418620 22420
rect 418488 22380 418494 22392
rect 418614 22380 418620 22392
rect 418672 22380 418678 22432
rect 217318 20000 217324 20052
rect 217376 20040 217382 20052
rect 371142 20040 371148 20052
rect 217376 20012 371148 20040
rect 217376 20000 217382 20012
rect 371142 20000 371148 20012
rect 371200 20000 371206 20052
rect 416314 19728 416320 19780
rect 416372 19768 416378 19780
rect 460658 19768 460664 19780
rect 416372 19740 460664 19768
rect 416372 19728 416378 19740
rect 460658 19728 460664 19740
rect 460716 19728 460722 19780
rect 405458 19660 405464 19712
rect 405516 19700 405522 19712
rect 488258 19700 488264 19712
rect 405516 19672 488264 19700
rect 405516 19660 405522 19672
rect 488258 19660 488264 19672
rect 488316 19660 488322 19712
rect 405090 19592 405096 19644
rect 405148 19632 405154 19644
rect 491018 19632 491024 19644
rect 405148 19604 491024 19632
rect 405148 19592 405154 19604
rect 491018 19592 491024 19604
rect 491076 19592 491082 19644
rect 405274 19524 405280 19576
rect 405332 19564 405338 19576
rect 493410 19564 493416 19576
rect 405332 19536 493416 19564
rect 405332 19524 405338 19536
rect 493410 19524 493416 19536
rect 493468 19524 493474 19576
rect 405550 19456 405556 19508
rect 405608 19496 405614 19508
rect 495894 19496 495900 19508
rect 405608 19468 495900 19496
rect 405608 19456 405614 19468
rect 495894 19456 495900 19468
rect 495952 19456 495958 19508
rect 17126 19388 17132 19440
rect 17184 19428 17190 19440
rect 52362 19428 52368 19440
rect 17184 19400 52368 19428
rect 17184 19388 17190 19400
rect 52362 19388 52368 19400
rect 52420 19388 52426 19440
rect 402698 19388 402704 19440
rect 402756 19428 402762 19440
rect 500954 19428 500960 19440
rect 402756 19400 500960 19428
rect 402756 19388 402762 19400
rect 500954 19388 500960 19400
rect 501012 19388 501018 19440
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 53466 19360 53472 19372
rect 15068 19332 53472 19360
rect 15068 19320 15074 19332
rect 53466 19320 53472 19332
rect 53524 19320 53530 19372
rect 188982 19320 188988 19372
rect 189040 19360 189046 19372
rect 285950 19360 285956 19372
rect 189040 19332 285956 19360
rect 189040 19320 189046 19332
rect 285950 19320 285956 19332
rect 286008 19320 286014 19372
rect 402790 19320 402796 19372
rect 402848 19360 402854 19372
rect 503530 19360 503536 19372
rect 402848 19332 503536 19360
rect 402848 19320 402854 19332
rect 503530 19320 503536 19332
rect 503588 19320 503594 19372
rect 103698 19252 103704 19304
rect 103756 19292 103762 19304
rect 176194 19292 176200 19304
rect 103756 19264 176200 19292
rect 103756 19252 103762 19264
rect 176194 19252 176200 19264
rect 176252 19252 176258 19304
rect 188798 19252 188804 19304
rect 188856 19292 188862 19304
rect 244274 19292 244280 19304
rect 188856 19264 244280 19292
rect 188856 19252 188862 19264
rect 244274 19252 244280 19264
rect 244332 19252 244338 19304
rect 415302 19252 415308 19304
rect 415360 19292 415366 19304
rect 447594 19292 447600 19304
rect 415360 19264 447600 19292
rect 415360 19252 415366 19264
rect 447594 19252 447600 19264
rect 447652 19252 447658 19304
rect 100938 19184 100944 19236
rect 100996 19224 101002 19236
rect 176286 19224 176292 19236
rect 100996 19196 176292 19224
rect 100996 19184 101002 19196
rect 176286 19184 176292 19196
rect 176344 19184 176350 19236
rect 190270 19184 190276 19236
rect 190328 19224 190334 19236
rect 246390 19224 246396 19236
rect 190328 19196 246396 19224
rect 190328 19184 190334 19196
rect 246390 19184 246396 19196
rect 246448 19184 246454 19236
rect 416222 19184 416228 19236
rect 416280 19224 416286 19236
rect 448698 19224 448704 19236
rect 416280 19196 448704 19224
rect 416280 19184 416286 19196
rect 448698 19184 448704 19196
rect 448756 19184 448762 19236
rect 95970 19116 95976 19168
rect 96028 19156 96034 19168
rect 176562 19156 176568 19168
rect 96028 19128 176568 19156
rect 96028 19116 96034 19128
rect 176562 19116 176568 19128
rect 176620 19116 176626 19168
rect 188522 19116 188528 19168
rect 188580 19156 188586 19168
rect 245286 19156 245292 19168
rect 188580 19128 245292 19156
rect 188580 19116 188586 19128
rect 245286 19116 245292 19128
rect 245344 19116 245350 19168
rect 416406 19116 416412 19168
rect 416464 19156 416470 19168
rect 455966 19156 455972 19168
rect 416464 19128 455972 19156
rect 416464 19116 416470 19128
rect 455966 19116 455972 19128
rect 456024 19116 456030 19168
rect 91002 19048 91008 19100
rect 91060 19088 91066 19100
rect 178586 19088 178592 19100
rect 91060 19060 178592 19088
rect 91060 19048 91066 19060
rect 178586 19048 178592 19060
rect 178644 19048 178650 19100
rect 188614 19048 188620 19100
rect 188672 19088 188678 19100
rect 248230 19088 248236 19100
rect 188672 19060 248236 19088
rect 188672 19048 188678 19060
rect 248230 19048 248236 19060
rect 248288 19048 248294 19100
rect 399478 19048 399484 19100
rect 399536 19088 399542 19100
rect 468294 19088 468300 19100
rect 399536 19060 468300 19088
rect 399536 19048 399542 19060
rect 468294 19048 468300 19060
rect 468352 19048 468358 19100
rect 86034 18980 86040 19032
rect 86092 19020 86098 19032
rect 179138 19020 179144 19032
rect 86092 18992 179144 19020
rect 86092 18980 86098 18992
rect 179138 18980 179144 18992
rect 179196 18980 179202 19032
rect 191742 18980 191748 19032
rect 191800 19020 191806 19032
rect 250070 19020 250076 19032
rect 191800 18992 250076 19020
rect 191800 18980 191806 18992
rect 250070 18980 250076 18992
rect 250128 18980 250134 19032
rect 399570 18980 399576 19032
rect 399628 19020 399634 19032
rect 470870 19020 470876 19032
rect 399628 18992 470876 19020
rect 399628 18980 399634 18992
rect 470870 18980 470876 18992
rect 470928 18980 470934 19032
rect 81066 18912 81072 18964
rect 81124 18952 81130 18964
rect 179322 18952 179328 18964
rect 81124 18924 179328 18952
rect 81124 18912 81130 18924
rect 179322 18912 179328 18924
rect 179380 18912 179386 18964
rect 187510 18912 187516 18964
rect 187568 18952 187574 18964
rect 247494 18952 247500 18964
rect 187568 18924 247500 18952
rect 187568 18912 187574 18924
rect 247494 18912 247500 18924
rect 247552 18912 247558 18964
rect 416038 18912 416044 18964
rect 416096 18952 416102 18964
rect 515766 18952 515772 18964
rect 416096 18924 515772 18952
rect 416096 18912 416102 18924
rect 515766 18912 515772 18924
rect 515824 18912 515830 18964
rect 76098 18844 76104 18896
rect 76156 18884 76162 18896
rect 179046 18884 179052 18896
rect 76156 18856 179052 18884
rect 76156 18844 76162 18856
rect 179046 18844 179052 18856
rect 179104 18844 179110 18896
rect 190178 18844 190184 18896
rect 190236 18884 190242 18896
rect 250622 18884 250628 18896
rect 190236 18856 250628 18884
rect 190236 18844 190242 18856
rect 250622 18844 250628 18856
rect 250680 18844 250686 18896
rect 402606 18844 402612 18896
rect 402664 18884 402670 18896
rect 505830 18884 505836 18896
rect 402664 18856 505836 18884
rect 402664 18844 402670 18856
rect 505830 18844 505836 18856
rect 505888 18844 505894 18896
rect 18414 18776 18420 18828
rect 18472 18816 18478 18828
rect 58158 18816 58164 18828
rect 18472 18788 58164 18816
rect 18472 18776 18478 18788
rect 58158 18776 58164 18788
rect 58216 18776 58222 18828
rect 73706 18776 73712 18828
rect 73764 18816 73770 18828
rect 181530 18816 181536 18828
rect 73764 18788 181536 18816
rect 73764 18776 73770 18788
rect 181530 18776 181536 18788
rect 181588 18776 181594 18828
rect 190362 18776 190368 18828
rect 190420 18816 190426 18828
rect 252278 18816 252284 18828
rect 190420 18788 252284 18816
rect 190420 18776 190426 18788
rect 252278 18776 252284 18788
rect 252336 18776 252342 18828
rect 402514 18776 402520 18828
rect 402572 18816 402578 18828
rect 508406 18816 508412 18828
rect 402572 18788 508412 18816
rect 402572 18776 402578 18788
rect 508406 18776 508412 18788
rect 508464 18776 508470 18828
rect 56042 18708 56048 18760
rect 56100 18748 56106 18760
rect 173618 18748 173624 18760
rect 56100 18720 173624 18748
rect 56100 18708 56106 18720
rect 173618 18708 173624 18720
rect 173676 18708 173682 18760
rect 191650 18708 191656 18760
rect 191708 18748 191714 18760
rect 253566 18748 253572 18760
rect 191708 18720 253572 18748
rect 191708 18708 191714 18720
rect 253566 18708 253572 18720
rect 253624 18708 253630 18760
rect 389910 18708 389916 18760
rect 389968 18748 389974 18760
rect 498470 18748 498476 18760
rect 389968 18720 498476 18748
rect 389968 18708 389974 18720
rect 498470 18708 498476 18720
rect 498528 18708 498534 18760
rect 53650 18640 53656 18692
rect 53708 18680 53714 18692
rect 173802 18680 173808 18692
rect 53708 18652 173808 18680
rect 53708 18640 53714 18652
rect 173802 18640 173808 18652
rect 173860 18640 173866 18692
rect 185854 18640 185860 18692
rect 185912 18680 185918 18692
rect 255958 18680 255964 18692
rect 185912 18652 255964 18680
rect 185912 18640 185918 18652
rect 255958 18640 255964 18652
rect 256016 18640 256022 18692
rect 389818 18640 389824 18692
rect 389876 18680 389882 18692
rect 523310 18680 523316 18692
rect 389876 18652 523316 18680
rect 389876 18640 389882 18652
rect 523310 18640 523316 18652
rect 523368 18640 523374 18692
rect 50890 18572 50896 18624
rect 50948 18612 50954 18624
rect 176378 18612 176384 18624
rect 50948 18584 176384 18612
rect 50948 18572 50954 18584
rect 176378 18572 176384 18584
rect 176436 18572 176442 18624
rect 185762 18572 185768 18624
rect 185820 18612 185826 18624
rect 258350 18612 258356 18624
rect 185820 18584 258356 18612
rect 185820 18572 185826 18584
rect 258350 18572 258356 18584
rect 258408 18572 258414 18624
rect 390002 18572 390008 18624
rect 390060 18612 390066 18624
rect 525886 18612 525892 18624
rect 390060 18584 525892 18612
rect 390060 18572 390066 18584
rect 525886 18572 525892 18584
rect 525944 18572 525950 18624
rect 106090 18504 106096 18556
rect 106148 18544 106154 18556
rect 176470 18544 176476 18556
rect 106148 18516 176476 18544
rect 106148 18504 106154 18516
rect 176470 18504 176476 18516
rect 176528 18504 176534 18556
rect 188706 18504 188712 18556
rect 188764 18544 188770 18556
rect 243078 18544 243084 18556
rect 188764 18516 243084 18544
rect 188764 18504 188770 18516
rect 243078 18504 243084 18516
rect 243136 18504 243142 18556
rect 418706 18504 418712 18556
rect 418764 18544 418770 18556
rect 450078 18544 450084 18556
rect 418764 18516 450084 18544
rect 418764 18504 418770 18516
rect 450078 18504 450084 18516
rect 450136 18504 450142 18556
rect 108666 18436 108672 18488
rect 108724 18476 108730 18488
rect 175918 18476 175924 18488
rect 108724 18448 175924 18476
rect 108724 18436 108730 18448
rect 175918 18436 175924 18448
rect 175976 18436 175982 18488
rect 188430 18436 188436 18488
rect 188488 18476 188494 18488
rect 235994 18476 236000 18488
rect 188488 18448 236000 18476
rect 188488 18436 188494 18448
rect 235994 18436 236000 18448
rect 236052 18436 236058 18488
rect 414566 18436 414572 18488
rect 414624 18476 414630 18488
rect 445662 18476 445668 18488
rect 414624 18448 445668 18476
rect 414624 18436 414630 18448
rect 445662 18436 445668 18448
rect 445720 18436 445726 18488
rect 113450 18368 113456 18420
rect 113508 18408 113514 18420
rect 176102 18408 176108 18420
rect 113508 18380 176108 18408
rect 113508 18368 113514 18380
rect 176102 18368 176108 18380
rect 176160 18368 176166 18420
rect 217410 18368 217416 18420
rect 217468 18408 217474 18420
rect 222194 18408 222200 18420
rect 217468 18380 222200 18408
rect 217468 18368 217474 18380
rect 222194 18368 222200 18380
rect 222252 18368 222258 18420
rect 415118 18368 415124 18420
rect 415176 18408 415182 18420
rect 444282 18408 444288 18420
rect 415176 18380 444288 18408
rect 415176 18368 415182 18380
rect 444282 18368 444288 18380
rect 444340 18368 444346 18420
rect 19058 17892 19064 17944
rect 19116 17932 19122 17944
rect 36538 17932 36544 17944
rect 19116 17904 36544 17932
rect 19116 17892 19122 17904
rect 36538 17892 36544 17904
rect 36596 17892 36602 17944
rect 62022 17892 62028 17944
rect 62080 17932 62086 17944
rect 173342 17932 173348 17944
rect 62080 17904 173348 17932
rect 62080 17892 62086 17904
rect 173342 17892 173348 17904
rect 173400 17892 173406 17944
rect 185670 17892 185676 17944
rect 185728 17932 185734 17944
rect 280154 17932 280160 17944
rect 185728 17904 280160 17932
rect 185728 17892 185734 17904
rect 280154 17892 280160 17904
rect 280212 17892 280218 17944
rect 402422 17892 402428 17944
rect 402480 17932 402486 17944
rect 458358 17932 458364 17944
rect 402480 17904 458364 17932
rect 402480 17892 402486 17904
rect 458358 17892 458364 17904
rect 458416 17892 458422 17944
rect 460658 17892 460664 17944
rect 460716 17932 460722 17944
rect 478874 17932 478880 17944
rect 460716 17904 478880 17932
rect 460716 17892 460722 17904
rect 478874 17892 478880 17904
rect 478932 17892 478938 17944
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 60458 17864 60464 17876
rect 19668 17836 60464 17864
rect 19668 17824 19674 17836
rect 60458 17824 60464 17836
rect 60516 17824 60522 17876
rect 64690 17824 64696 17876
rect 64748 17864 64754 17876
rect 173434 17864 173440 17876
rect 64748 17836 173440 17864
rect 64748 17824 64754 17836
rect 173434 17824 173440 17836
rect 173492 17824 173498 17876
rect 187602 17824 187608 17876
rect 187660 17864 187666 17876
rect 277394 17864 277400 17876
rect 187660 17836 277400 17864
rect 187660 17824 187666 17836
rect 277394 17824 277400 17836
rect 277452 17824 277458 17876
rect 444282 17824 444288 17876
rect 444340 17864 444346 17876
rect 462314 17864 462320 17876
rect 444340 17836 462320 17864
rect 444340 17824 444346 17836
rect 462314 17824 462320 17836
rect 462372 17824 462378 17876
rect 18506 17756 18512 17808
rect 18564 17796 18570 17808
rect 55950 17796 55956 17808
rect 18564 17768 55956 17796
rect 18564 17756 18570 17768
rect 55950 17756 55956 17768
rect 56008 17796 56014 17808
rect 56502 17796 56508 17808
rect 56008 17768 56508 17796
rect 56008 17756 56014 17768
rect 56502 17756 56508 17768
rect 56560 17756 56566 17808
rect 66162 17756 66168 17808
rect 66220 17796 66226 17808
rect 173158 17796 173164 17808
rect 66220 17768 173164 17796
rect 66220 17756 66226 17768
rect 173158 17756 173164 17768
rect 173216 17756 173222 17808
rect 191466 17756 191472 17808
rect 191524 17796 191530 17808
rect 273254 17796 273260 17808
rect 191524 17768 273260 17796
rect 191524 17756 191530 17768
rect 273254 17756 273260 17768
rect 273312 17756 273318 17808
rect 410518 17756 410524 17808
rect 410576 17796 410582 17808
rect 455414 17796 455420 17808
rect 410576 17768 455420 17796
rect 410576 17756 410582 17768
rect 455414 17756 455420 17768
rect 455472 17756 455478 17808
rect 455966 17756 455972 17808
rect 456024 17796 456030 17808
rect 473354 17796 473360 17808
rect 456024 17768 473360 17796
rect 456024 17756 456030 17768
rect 473354 17756 473360 17768
rect 473412 17756 473418 17808
rect 18598 17688 18604 17740
rect 18656 17728 18662 17740
rect 53834 17728 53840 17740
rect 18656 17700 53840 17728
rect 18656 17688 18662 17700
rect 53834 17688 53840 17700
rect 53892 17688 53898 17740
rect 68922 17688 68928 17740
rect 68980 17728 68986 17740
rect 173250 17728 173256 17740
rect 68980 17700 173256 17728
rect 68980 17688 68986 17700
rect 173250 17688 173256 17700
rect 173308 17688 173314 17740
rect 183462 17688 183468 17740
rect 183520 17728 183526 17740
rect 264974 17728 264980 17740
rect 183520 17700 264980 17728
rect 183520 17688 183526 17700
rect 264974 17688 264980 17700
rect 265032 17688 265038 17740
rect 414474 17688 414480 17740
rect 414532 17728 414538 17740
rect 456794 17728 456800 17740
rect 414532 17700 456800 17728
rect 414532 17688 414538 17700
rect 456794 17688 456800 17700
rect 456852 17688 456858 17740
rect 16206 17620 16212 17672
rect 16264 17660 16270 17672
rect 51442 17660 51448 17672
rect 16264 17632 51448 17660
rect 16264 17620 16270 17632
rect 51442 17620 51448 17632
rect 51500 17620 51506 17672
rect 78582 17620 78588 17672
rect 78640 17660 78646 17672
rect 178770 17660 178776 17672
rect 78640 17632 178776 17660
rect 78640 17620 78646 17632
rect 178770 17620 178776 17632
rect 178828 17620 178834 17672
rect 183370 17620 183376 17672
rect 183428 17660 183434 17672
rect 263594 17660 263600 17672
rect 183428 17632 263600 17660
rect 183428 17620 183434 17632
rect 263594 17620 263600 17632
rect 263652 17620 263658 17672
rect 445662 17620 445668 17672
rect 445720 17660 445726 17672
rect 463694 17660 463700 17672
rect 445720 17632 463700 17660
rect 445720 17620 445726 17632
rect 463694 17620 463700 17632
rect 463752 17620 463758 17672
rect 16390 17552 16396 17604
rect 16448 17592 16454 17604
rect 48682 17592 48688 17604
rect 16448 17564 48688 17592
rect 16448 17552 16454 17564
rect 48682 17552 48688 17564
rect 48740 17592 48746 17604
rect 49602 17592 49608 17604
rect 48740 17564 49608 17592
rect 48740 17552 48746 17564
rect 49602 17552 49608 17564
rect 49660 17552 49666 17604
rect 53466 17552 53472 17604
rect 53524 17592 53530 17604
rect 71774 17592 71780 17604
rect 53524 17564 71780 17592
rect 53524 17552 53530 17564
rect 71774 17552 71780 17564
rect 71832 17552 71838 17604
rect 191834 17552 191840 17604
rect 191892 17592 191898 17604
rect 270494 17592 270500 17604
rect 191892 17564 270500 17592
rect 191892 17552 191898 17564
rect 270494 17552 270500 17564
rect 270552 17552 270558 17604
rect 448698 17552 448704 17604
rect 448756 17592 448762 17604
rect 466454 17592 466460 17604
rect 448756 17564 466460 17592
rect 448756 17552 448762 17564
rect 466454 17552 466460 17564
rect 466512 17552 466518 17604
rect 15102 17484 15108 17536
rect 15160 17524 15166 17536
rect 47578 17524 47584 17536
rect 15160 17496 47584 17524
rect 15160 17484 15166 17496
rect 47578 17484 47584 17496
rect 47636 17524 47642 17536
rect 48222 17524 48228 17536
rect 47636 17496 48228 17524
rect 47636 17484 47642 17496
rect 48222 17484 48228 17496
rect 48280 17484 48286 17536
rect 50154 17484 50160 17536
rect 50212 17524 50218 17536
rect 67634 17524 67640 17536
rect 50212 17496 67640 17524
rect 50212 17484 50218 17496
rect 67634 17484 67640 17496
rect 67692 17484 67698 17536
rect 83826 17484 83832 17536
rect 83884 17524 83890 17536
rect 178678 17524 178684 17536
rect 83884 17496 178684 17524
rect 83884 17484 83890 17496
rect 178678 17484 178684 17496
rect 178736 17484 178742 17536
rect 185946 17484 185952 17536
rect 186004 17524 186010 17536
rect 260834 17524 260840 17536
rect 186004 17496 260840 17524
rect 186004 17484 186010 17496
rect 260834 17484 260840 17496
rect 260892 17484 260898 17536
rect 419258 17484 419264 17536
rect 419316 17524 419322 17536
rect 443086 17524 443092 17536
rect 419316 17496 443092 17524
rect 419316 17484 419322 17496
rect 443086 17484 443092 17496
rect 443144 17524 443150 17536
rect 443144 17496 444880 17524
rect 443144 17484 443150 17496
rect 19242 17416 19248 17468
rect 19300 17456 19306 17468
rect 50172 17456 50200 17484
rect 19300 17428 50200 17456
rect 19300 17416 19306 17428
rect 60458 17416 60464 17468
rect 60516 17456 60522 17468
rect 78674 17456 78680 17468
rect 60516 17428 78680 17456
rect 60516 17416 60522 17428
rect 78674 17416 78680 17428
rect 78732 17416 78738 17468
rect 88242 17416 88248 17468
rect 88300 17456 88306 17468
rect 178862 17456 178868 17468
rect 88300 17428 178868 17456
rect 88300 17416 88306 17428
rect 178862 17416 178868 17428
rect 178920 17416 178926 17468
rect 184750 17416 184756 17468
rect 184808 17456 184814 17468
rect 259546 17456 259552 17468
rect 184808 17428 259552 17456
rect 184808 17416 184814 17428
rect 259546 17416 259552 17428
rect 259604 17416 259610 17468
rect 417050 17416 417056 17468
rect 417108 17456 417114 17468
rect 441706 17456 441712 17468
rect 417108 17428 441712 17456
rect 417108 17416 417114 17428
rect 441706 17416 441712 17428
rect 441764 17416 441770 17468
rect 19426 17348 19432 17400
rect 19484 17388 19490 17400
rect 19484 17360 45554 17388
rect 19484 17348 19490 17360
rect 18322 17280 18328 17332
rect 18380 17320 18386 17332
rect 18380 17292 42288 17320
rect 18380 17280 18386 17292
rect 19518 17212 19524 17264
rect 19576 17252 19582 17264
rect 19576 17224 41920 17252
rect 19576 17212 19582 17224
rect 19702 17144 19708 17196
rect 19760 17184 19766 17196
rect 19760 17156 41460 17184
rect 19760 17144 19766 17156
rect 18874 17076 18880 17128
rect 18932 17116 18938 17128
rect 38654 17116 38660 17128
rect 18932 17088 38660 17116
rect 18932 17076 18938 17088
rect 38654 17076 38660 17088
rect 38712 17076 38718 17128
rect 41432 17048 41460 17156
rect 41892 17116 41920 17224
rect 42260 17184 42288 17292
rect 45526 17252 45554 17360
rect 49602 17348 49608 17400
rect 49660 17388 49666 17400
rect 67634 17388 67640 17400
rect 49660 17360 67640 17388
rect 49660 17348 49666 17360
rect 67634 17348 67640 17360
rect 67692 17348 67698 17400
rect 69658 17348 69664 17400
rect 69716 17388 69722 17400
rect 75914 17388 75920 17400
rect 69716 17360 75920 17388
rect 69716 17348 69722 17360
rect 75914 17348 75920 17360
rect 75972 17348 75978 17400
rect 93578 17348 93584 17400
rect 93636 17388 93642 17400
rect 178954 17388 178960 17400
rect 93636 17360 178960 17388
rect 93636 17348 93642 17360
rect 178954 17348 178960 17360
rect 179012 17348 179018 17400
rect 186038 17348 186044 17400
rect 186096 17388 186102 17400
rect 259454 17388 259460 17400
rect 186096 17360 259460 17388
rect 186096 17348 186102 17360
rect 259454 17348 259460 17360
rect 259512 17348 259518 17400
rect 418062 17348 418068 17400
rect 418120 17388 418126 17400
rect 440234 17388 440240 17400
rect 418120 17360 440240 17388
rect 418120 17348 418126 17360
rect 440234 17348 440240 17360
rect 440292 17348 440298 17400
rect 444852 17388 444880 17496
rect 450078 17484 450084 17536
rect 450136 17524 450142 17536
rect 467834 17524 467840 17536
rect 450136 17496 467840 17524
rect 450136 17484 450142 17496
rect 467834 17484 467840 17496
rect 467892 17484 467898 17536
rect 447594 17416 447600 17468
rect 447652 17456 447658 17468
rect 465074 17456 465080 17468
rect 447652 17428 465080 17456
rect 447652 17416 447658 17428
rect 465074 17416 465080 17428
rect 465132 17416 465138 17468
rect 459462 17388 459468 17400
rect 444852 17360 459468 17388
rect 459462 17348 459468 17360
rect 459520 17348 459526 17400
rect 48222 17280 48228 17332
rect 48280 17320 48286 17332
rect 66254 17320 66260 17332
rect 48280 17292 66260 17320
rect 48280 17280 48286 17292
rect 66254 17280 66260 17292
rect 66312 17280 66318 17332
rect 99282 17280 99288 17332
rect 99340 17320 99346 17332
rect 176010 17320 176016 17332
rect 99340 17292 176016 17320
rect 99340 17280 99346 17292
rect 176010 17280 176016 17292
rect 176068 17280 176074 17332
rect 186130 17280 186136 17332
rect 186188 17320 186194 17332
rect 258074 17320 258080 17332
rect 186188 17292 258080 17320
rect 186188 17280 186194 17292
rect 258074 17280 258080 17292
rect 258132 17280 258138 17332
rect 419718 17280 419724 17332
rect 419776 17320 419782 17332
rect 438854 17320 438860 17332
rect 419776 17292 438860 17320
rect 419776 17280 419782 17292
rect 438854 17280 438860 17292
rect 438912 17280 438918 17332
rect 456794 17280 456800 17332
rect 456852 17320 456858 17332
rect 458082 17320 458088 17332
rect 456852 17292 458088 17320
rect 456852 17280 456858 17292
rect 458082 17280 458088 17292
rect 458140 17320 458146 17332
rect 476114 17320 476120 17332
rect 458140 17292 476120 17320
rect 458140 17280 458146 17292
rect 476114 17280 476120 17292
rect 476172 17280 476178 17332
rect 46658 17252 46664 17264
rect 45526 17224 46664 17252
rect 46658 17212 46664 17224
rect 46716 17252 46722 17264
rect 65058 17252 65064 17264
rect 46716 17224 65064 17252
rect 46716 17212 46722 17224
rect 65058 17212 65064 17224
rect 65116 17212 65122 17264
rect 111702 17212 111708 17264
rect 111760 17252 111766 17264
rect 157978 17252 157984 17264
rect 111760 17224 157984 17252
rect 111760 17212 111766 17224
rect 157978 17212 157984 17224
rect 158036 17212 158042 17264
rect 184842 17212 184848 17264
rect 184900 17252 184906 17264
rect 256694 17252 256700 17264
rect 184900 17224 256700 17252
rect 184900 17212 184906 17224
rect 256694 17212 256700 17224
rect 256752 17212 256758 17264
rect 419810 17212 419816 17264
rect 419868 17252 419874 17264
rect 437474 17252 437480 17264
rect 419868 17224 437480 17252
rect 419868 17212 419874 17224
rect 437474 17212 437480 17224
rect 437532 17212 437538 17264
rect 465074 17252 465080 17264
rect 451246 17224 465080 17252
rect 45370 17184 45376 17196
rect 42260 17156 45376 17184
rect 45370 17144 45376 17156
rect 45428 17184 45434 17196
rect 63494 17184 63500 17196
rect 45428 17156 63500 17184
rect 45428 17144 45434 17156
rect 63494 17144 63500 17156
rect 63552 17144 63558 17196
rect 71682 17144 71688 17196
rect 71740 17184 71746 17196
rect 170398 17184 170404 17196
rect 71740 17156 170404 17184
rect 71740 17144 71746 17156
rect 170398 17144 170404 17156
rect 170456 17144 170462 17196
rect 186222 17144 186228 17196
rect 186280 17184 186286 17196
rect 255314 17184 255320 17196
rect 186280 17156 255320 17184
rect 186280 17144 186286 17156
rect 255314 17144 255320 17156
rect 255372 17144 255378 17196
rect 419166 17144 419172 17196
rect 419224 17184 419230 17196
rect 436094 17184 436100 17196
rect 419224 17156 436100 17184
rect 419224 17144 419230 17156
rect 436094 17144 436100 17156
rect 436152 17144 436158 17196
rect 44174 17116 44180 17128
rect 41892 17088 44180 17116
rect 44174 17076 44180 17088
rect 44232 17116 44238 17128
rect 62114 17116 62120 17128
rect 44232 17088 62120 17116
rect 44232 17076 44238 17088
rect 62114 17076 62120 17088
rect 62172 17076 62178 17128
rect 218698 17076 218704 17128
rect 218756 17116 218762 17128
rect 282914 17116 282920 17128
rect 218756 17088 282920 17116
rect 218756 17076 218762 17088
rect 282914 17076 282920 17088
rect 282972 17076 282978 17128
rect 418982 17076 418988 17128
rect 419040 17116 419046 17128
rect 436278 17116 436284 17128
rect 419040 17088 436284 17116
rect 419040 17076 419046 17088
rect 436278 17076 436284 17088
rect 436336 17076 436342 17128
rect 43070 17048 43076 17060
rect 41432 17020 43076 17048
rect 43070 17008 43076 17020
rect 43128 17048 43134 17060
rect 60734 17048 60740 17060
rect 43128 17020 60740 17048
rect 43128 17008 43134 17020
rect 60734 17008 60740 17020
rect 60792 17008 60798 17060
rect 191098 17008 191104 17060
rect 191156 17048 191162 17060
rect 251174 17048 251180 17060
rect 191156 17020 251180 17048
rect 191156 17008 191162 17020
rect 251174 17008 251180 17020
rect 251232 17008 251238 17060
rect 393958 17008 393964 17060
rect 394016 17048 394022 17060
rect 447134 17048 447140 17060
rect 394016 17020 447140 17048
rect 394016 17008 394022 17020
rect 447134 17008 447140 17020
rect 447192 17008 447198 17060
rect 51442 16940 51448 16992
rect 51500 16980 51506 16992
rect 69014 16980 69020 16992
rect 51500 16952 69020 16980
rect 51500 16940 51506 16952
rect 69014 16940 69020 16952
rect 69072 16940 69078 16992
rect 414382 16940 414388 16992
rect 414440 16980 414446 16992
rect 446490 16980 446496 16992
rect 414440 16952 446496 16980
rect 414440 16940 414446 16952
rect 446490 16940 446496 16952
rect 446548 16980 446554 16992
rect 451246 16980 451274 17224
rect 465074 17212 465080 17224
rect 465132 17212 465138 17264
rect 469306 16980 469312 16992
rect 446548 16952 451274 16980
rect 460906 16952 469312 16980
rect 446548 16940 446554 16952
rect 16482 16872 16488 16924
rect 16540 16912 16546 16924
rect 59538 16912 59544 16924
rect 16540 16884 59544 16912
rect 16540 16872 16546 16884
rect 59538 16872 59544 16884
rect 59596 16912 59602 16924
rect 77294 16912 77300 16924
rect 59596 16884 77300 16912
rect 59596 16872 59602 16884
rect 77294 16872 77300 16884
rect 77352 16872 77358 16924
rect 418430 16872 418436 16924
rect 418488 16912 418494 16924
rect 449894 16912 449900 16924
rect 418488 16884 449900 16912
rect 418488 16872 418494 16884
rect 449894 16872 449900 16884
rect 449952 16872 449958 16924
rect 451274 16872 451280 16924
rect 451332 16912 451338 16924
rect 460906 16912 460934 16952
rect 469306 16940 469312 16952
rect 469364 16940 469370 16992
rect 451332 16884 460934 16912
rect 451332 16872 451338 16884
rect 469214 16872 469220 16924
rect 469272 16912 469278 16924
rect 473446 16912 473452 16924
rect 469272 16884 473452 16912
rect 469272 16872 469278 16884
rect 473446 16872 473452 16884
rect 473504 16872 473510 16924
rect 56502 16804 56508 16856
rect 56560 16844 56566 16856
rect 73154 16844 73160 16856
rect 56560 16816 73160 16844
rect 56560 16804 56566 16816
rect 73154 16804 73160 16816
rect 73212 16804 73218 16856
rect 457346 16804 457352 16856
rect 457404 16844 457410 16856
rect 474734 16844 474740 16856
rect 457404 16816 474740 16844
rect 457404 16804 457410 16816
rect 474734 16804 474740 16816
rect 474792 16804 474798 16856
rect 57882 16736 57888 16788
rect 57940 16776 57946 16788
rect 74810 16776 74816 16788
rect 57940 16748 74816 16776
rect 57940 16736 57946 16748
rect 74810 16736 74816 16748
rect 74868 16736 74874 16788
rect 451366 16736 451372 16788
rect 451424 16776 451430 16788
rect 452286 16776 452292 16788
rect 451424 16748 452292 16776
rect 451424 16736 451430 16748
rect 452286 16736 452292 16748
rect 452344 16776 452350 16788
rect 470870 16776 470876 16788
rect 452344 16748 470876 16776
rect 452344 16736 452350 16748
rect 470870 16736 470876 16748
rect 470928 16736 470934 16788
rect 52362 16668 52368 16720
rect 52420 16708 52426 16720
rect 70394 16708 70400 16720
rect 52420 16680 70400 16708
rect 52420 16668 52426 16680
rect 70394 16668 70400 16680
rect 70452 16668 70458 16720
rect 452654 16668 452660 16720
rect 452712 16708 452718 16720
rect 453482 16708 453488 16720
rect 452712 16680 453488 16708
rect 452712 16668 452718 16680
rect 453482 16668 453488 16680
rect 453540 16708 453546 16720
rect 471974 16708 471980 16720
rect 453540 16680 471980 16708
rect 453540 16668 453546 16680
rect 471974 16668 471980 16680
rect 472032 16668 472038 16720
rect 477494 16640 477500 16652
rect 458652 16612 477500 16640
rect 125962 16532 125968 16584
rect 126020 16572 126026 16584
rect 388070 16572 388076 16584
rect 126020 16544 388076 16572
rect 126020 16532 126026 16544
rect 388070 16532 388076 16544
rect 388128 16532 388134 16584
rect 416130 16532 416136 16584
rect 416188 16572 416194 16584
rect 458266 16572 458272 16584
rect 416188 16544 458272 16572
rect 416188 16532 416194 16544
rect 458266 16532 458272 16544
rect 458324 16572 458330 16584
rect 458652 16572 458680 16612
rect 477494 16600 477500 16612
rect 477552 16600 477558 16652
rect 458324 16544 458680 16572
rect 458324 16532 458330 16544
rect 418338 16464 418344 16516
rect 418396 16504 418402 16516
rect 457346 16504 457352 16516
rect 418396 16476 457352 16504
rect 418396 16464 418402 16476
rect 457346 16464 457352 16476
rect 457404 16464 457410 16516
rect 419902 16396 419908 16448
rect 419960 16436 419966 16448
rect 454034 16436 454040 16448
rect 419960 16408 454040 16436
rect 419960 16396 419966 16408
rect 454034 16396 454040 16408
rect 454092 16436 454098 16448
rect 469214 16436 469220 16448
rect 454092 16408 469220 16436
rect 454092 16396 454098 16408
rect 469214 16396 469220 16408
rect 469272 16396 469278 16448
rect 417970 16328 417976 16380
rect 418028 16368 418034 16380
rect 451274 16368 451280 16380
rect 418028 16340 451280 16368
rect 418028 16328 418034 16340
rect 451274 16328 451280 16340
rect 451332 16328 451338 16380
rect 419994 16260 420000 16312
rect 420052 16300 420058 16312
rect 452654 16300 452660 16312
rect 420052 16272 452660 16300
rect 420052 16260 420058 16272
rect 452654 16260 452660 16272
rect 452712 16260 452718 16312
rect 418614 16192 418620 16244
rect 418672 16232 418678 16244
rect 451366 16232 451372 16244
rect 418672 16204 451372 16232
rect 418672 16192 418678 16204
rect 451366 16192 451372 16204
rect 451424 16192 451430 16244
rect 359550 15920 359556 15972
rect 359608 15960 359614 15972
rect 420914 15960 420920 15972
rect 359608 15932 420920 15960
rect 359608 15920 359614 15932
rect 420914 15920 420920 15932
rect 420972 15920 420978 15972
rect 130562 15852 130568 15904
rect 130620 15892 130626 15904
rect 198734 15892 198740 15904
rect 130620 15864 198740 15892
rect 130620 15852 130626 15864
rect 198734 15852 198740 15864
rect 198792 15852 198798 15904
rect 363598 15852 363604 15904
rect 363656 15892 363662 15904
rect 432046 15892 432052 15904
rect 363656 15864 432052 15892
rect 363656 15852 363662 15864
rect 432046 15852 432052 15864
rect 432104 15852 432110 15904
rect 358354 14492 358360 14544
rect 358412 14532 358418 14544
rect 423674 14532 423680 14544
rect 358412 14504 423680 14532
rect 358412 14492 358418 14504
rect 423674 14492 423680 14504
rect 423732 14492 423738 14544
rect 126974 14424 126980 14476
rect 127032 14464 127038 14476
rect 197446 14464 197452 14476
rect 127032 14436 197452 14464
rect 127032 14424 127038 14436
rect 197446 14424 197452 14436
rect 197504 14424 197510 14476
rect 358170 14424 358176 14476
rect 358228 14464 358234 14476
rect 442626 14464 442632 14476
rect 358228 14436 442632 14464
rect 358228 14424 358234 14436
rect 442626 14424 442632 14436
rect 442684 14424 442690 14476
rect 362954 13064 362960 13116
rect 363012 13104 363018 13116
rect 552658 13104 552664 13116
rect 363012 13076 552664 13104
rect 363012 13064 363018 13076
rect 552658 13064 552664 13076
rect 552716 13064 552722 13116
rect 357434 11840 357440 11892
rect 357492 11880 357498 11892
rect 357492 11852 357664 11880
rect 357492 11840 357498 11852
rect 357636 11552 357664 11852
rect 360930 11772 360936 11824
rect 360988 11812 360994 11824
rect 428458 11812 428464 11824
rect 360988 11784 428464 11812
rect 360988 11772 360994 11784
rect 428458 11772 428464 11784
rect 428516 11772 428522 11824
rect 359458 11704 359464 11756
rect 359516 11744 359522 11756
rect 470594 11744 470600 11756
rect 359516 11716 470600 11744
rect 359516 11704 359522 11716
rect 470594 11704 470600 11716
rect 470652 11704 470658 11756
rect 357618 11500 357624 11552
rect 357676 11500 357682 11552
rect 128170 10276 128176 10328
rect 128228 10316 128234 10328
rect 195238 10316 195244 10328
rect 128228 10288 195244 10316
rect 128228 10276 128234 10288
rect 195238 10276 195244 10288
rect 195296 10276 195302 10328
rect 361574 10276 361580 10328
rect 361632 10316 361638 10328
rect 548610 10316 548616 10328
rect 361632 10288 548616 10316
rect 361632 10276 361638 10288
rect 548610 10276 548616 10288
rect 548668 10276 548674 10328
rect 360194 8916 360200 8968
rect 360252 8956 360258 8968
rect 545482 8956 545488 8968
rect 360252 8928 545488 8956
rect 360252 8916 360258 8928
rect 545482 8916 545488 8928
rect 545540 8916 545546 8968
rect 218882 8304 218888 8356
rect 218940 8344 218946 8356
rect 219066 8344 219072 8356
rect 218940 8316 219072 8344
rect 218940 8304 218946 8316
rect 219066 8304 219072 8316
rect 219124 8304 219130 8356
rect 357158 7624 357164 7676
rect 357216 7664 357222 7676
rect 527818 7664 527824 7676
rect 357216 7636 527824 7664
rect 357216 7624 357222 7636
rect 527818 7624 527824 7636
rect 527876 7624 527882 7676
rect 158898 7556 158904 7608
rect 158956 7596 158962 7608
rect 209774 7596 209780 7608
rect 158956 7568 209780 7596
rect 158956 7556 158962 7568
rect 209774 7556 209780 7568
rect 209832 7556 209838 7608
rect 218054 7556 218060 7608
rect 218112 7596 218118 7608
rect 219250 7596 219256 7608
rect 218112 7568 219256 7596
rect 218112 7556 218118 7568
rect 219250 7556 219256 7568
rect 219308 7556 219314 7608
rect 356974 7556 356980 7608
rect 357032 7596 357038 7608
rect 531314 7596 531320 7608
rect 357032 7568 531320 7596
rect 357032 7556 357038 7568
rect 531314 7556 531320 7568
rect 531372 7556 531378 7608
rect 216214 6332 216220 6384
rect 216272 6372 216278 6384
rect 293678 6372 293684 6384
rect 216272 6344 293684 6372
rect 216272 6332 216278 6344
rect 293678 6332 293684 6344
rect 293736 6332 293742 6384
rect 219710 6264 219716 6316
rect 219768 6304 219774 6316
rect 300762 6304 300768 6316
rect 219768 6276 300768 6304
rect 219768 6264 219774 6276
rect 300762 6264 300768 6276
rect 300820 6264 300826 6316
rect 216306 6196 216312 6248
rect 216364 6236 216370 6248
rect 297266 6236 297272 6248
rect 216364 6208 297272 6236
rect 216364 6196 216370 6208
rect 297266 6196 297272 6208
rect 297324 6196 297330 6248
rect 411990 6196 411996 6248
rect 412048 6236 412054 6248
rect 524230 6236 524236 6248
rect 412048 6208 524236 6236
rect 412048 6196 412054 6208
rect 524230 6196 524236 6208
rect 524288 6196 524294 6248
rect 169570 6128 169576 6180
rect 169628 6168 169634 6180
rect 213914 6168 213920 6180
rect 169628 6140 213920 6168
rect 169628 6128 169634 6140
rect 213914 6128 213920 6140
rect 213972 6128 213978 6180
rect 218974 6128 218980 6180
rect 219032 6168 219038 6180
rect 304350 6168 304356 6180
rect 219032 6140 304356 6168
rect 219032 6128 219038 6140
rect 304350 6128 304356 6140
rect 304408 6128 304414 6180
rect 357618 6128 357624 6180
rect 357676 6168 357682 6180
rect 538398 6168 538404 6180
rect 357676 6140 538404 6168
rect 357676 6128 357682 6140
rect 538398 6128 538404 6140
rect 538456 6128 538462 6180
rect 356698 5244 356704 5296
rect 356756 5284 356762 5296
rect 488810 5284 488816 5296
rect 356756 5256 488816 5284
rect 356756 5244 356762 5256
rect 488810 5244 488816 5256
rect 488868 5244 488874 5296
rect 360838 5176 360844 5228
rect 360896 5216 360902 5228
rect 495894 5216 495900 5228
rect 360896 5188 495900 5216
rect 360896 5176 360902 5188
rect 495894 5176 495900 5188
rect 495952 5176 495958 5228
rect 356790 5108 356796 5160
rect 356848 5148 356854 5160
rect 502978 5148 502984 5160
rect 356848 5120 502984 5148
rect 356848 5108 356854 5120
rect 502978 5108 502984 5120
rect 503036 5108 503042 5160
rect 358262 5040 358268 5092
rect 358320 5080 358326 5092
rect 506474 5080 506480 5092
rect 358320 5052 506480 5080
rect 358320 5040 358326 5052
rect 506474 5040 506480 5052
rect 506532 5040 506538 5092
rect 358078 4972 358084 5024
rect 358136 5012 358142 5024
rect 513558 5012 513564 5024
rect 358136 4984 513564 5012
rect 358136 4972 358142 4984
rect 513558 4972 513564 4984
rect 513616 4972 513622 5024
rect 364334 4904 364340 4956
rect 364392 4944 364398 4956
rect 556154 4944 556160 4956
rect 364392 4916 556160 4944
rect 364392 4904 364398 4916
rect 556154 4904 556160 4916
rect 556212 4904 556218 4956
rect 365714 4836 365720 4888
rect 365772 4876 365778 4888
rect 559742 4876 559748 4888
rect 365772 4848 559748 4876
rect 365772 4836 365778 4848
rect 559742 4836 559748 4848
rect 559800 4836 559806 4888
rect 125870 4768 125876 4820
rect 125928 4808 125934 4820
rect 194594 4808 194600 4820
rect 125928 4780 194600 4808
rect 125928 4768 125934 4780
rect 194594 4768 194600 4780
rect 194652 4768 194658 4820
rect 563238 4808 563244 4820
rect 373966 4780 563244 4808
rect 367094 4700 367100 4752
rect 367152 4740 367158 4752
rect 373966 4740 373994 4780
rect 563238 4768 563244 4780
rect 563296 4768 563302 4820
rect 367152 4712 373994 4740
rect 367152 4700 367158 4712
rect 217962 4088 217968 4140
rect 218020 4128 218026 4140
rect 237006 4128 237012 4140
rect 218020 4100 237012 4128
rect 218020 4088 218026 4100
rect 237006 4088 237012 4100
rect 237064 4088 237070 4140
rect 343358 4088 343364 4140
rect 343416 4128 343422 4140
rect 359182 4128 359188 4140
rect 343416 4100 359188 4128
rect 343416 4088 343422 4100
rect 359182 4088 359188 4100
rect 359240 4088 359246 4140
rect 414658 4088 414664 4140
rect 414716 4128 414722 4140
rect 449802 4128 449808 4140
rect 414716 4100 449808 4128
rect 414716 4088 414722 4100
rect 449802 4088 449808 4100
rect 449860 4088 449866 4140
rect 217870 4020 217876 4072
rect 217928 4060 217934 4072
rect 240502 4060 240508 4072
rect 217928 4032 240508 4060
rect 217928 4020 217934 4032
rect 240502 4020 240508 4032
rect 240560 4020 240566 4072
rect 339862 4020 339868 4072
rect 339920 4060 339926 4072
rect 357066 4060 357072 4072
rect 339920 4032 357072 4060
rect 339920 4020 339926 4032
rect 357066 4020 357072 4032
rect 357124 4020 357130 4072
rect 416590 4020 416596 4072
rect 416648 4060 416654 4072
rect 453298 4060 453304 4072
rect 416648 4032 453304 4060
rect 416648 4020 416654 4032
rect 453298 4020 453304 4032
rect 453356 4020 453362 4072
rect 217778 3952 217784 4004
rect 217836 3992 217842 4004
rect 244090 3992 244096 4004
rect 217836 3964 244096 3992
rect 217836 3952 217842 3964
rect 244090 3952 244096 3964
rect 244148 3952 244154 4004
rect 336274 3952 336280 4004
rect 336332 3992 336338 4004
rect 357894 3992 357900 4004
rect 336332 3964 357900 3992
rect 336332 3952 336338 3964
rect 357894 3952 357900 3964
rect 357952 3952 357958 4004
rect 411898 3952 411904 4004
rect 411956 3992 411962 4004
rect 456886 3992 456892 4004
rect 411956 3964 456892 3992
rect 411956 3952 411962 3964
rect 456886 3952 456892 3964
rect 456944 3952 456950 4004
rect 217686 3884 217692 3936
rect 217744 3924 217750 3936
rect 247586 3924 247592 3936
rect 217744 3896 247592 3924
rect 217744 3884 217750 3896
rect 247586 3884 247592 3896
rect 247644 3884 247650 3936
rect 332686 3884 332692 3936
rect 332744 3924 332750 3936
rect 357710 3924 357716 3936
rect 332744 3896 357716 3924
rect 332744 3884 332750 3896
rect 357710 3884 357716 3896
rect 357768 3884 357774 3936
rect 413830 3884 413836 3936
rect 413888 3924 413894 3936
rect 460382 3924 460388 3936
rect 413888 3896 460388 3924
rect 413888 3884 413894 3896
rect 460382 3884 460388 3896
rect 460440 3884 460446 3936
rect 155402 3816 155408 3868
rect 155460 3856 155466 3868
rect 175826 3856 175832 3868
rect 155460 3828 175832 3856
rect 155460 3816 155466 3828
rect 175826 3816 175832 3828
rect 175884 3816 175890 3868
rect 219342 3816 219348 3868
rect 219400 3856 219406 3868
rect 251174 3856 251180 3868
rect 219400 3828 251180 3856
rect 219400 3816 219406 3828
rect 251174 3816 251180 3828
rect 251232 3816 251238 3868
rect 329190 3816 329196 3868
rect 329248 3856 329254 3868
rect 357434 3856 357440 3868
rect 329248 3828 357440 3856
rect 329248 3816 329254 3828
rect 357434 3816 357440 3828
rect 357492 3816 357498 3868
rect 418798 3816 418804 3868
rect 418856 3856 418862 3868
rect 467466 3856 467472 3868
rect 418856 3828 467472 3856
rect 418856 3816 418862 3828
rect 467466 3816 467472 3828
rect 467524 3816 467530 3868
rect 151814 3748 151820 3800
rect 151872 3788 151878 3800
rect 174538 3788 174544 3800
rect 151872 3760 174544 3788
rect 151872 3748 151878 3760
rect 174538 3748 174544 3760
rect 174596 3748 174602 3800
rect 215202 3748 215208 3800
rect 215260 3788 215266 3800
rect 254670 3788 254676 3800
rect 215260 3760 254676 3788
rect 215260 3748 215266 3760
rect 254670 3748 254676 3760
rect 254728 3748 254734 3800
rect 325602 3748 325608 3800
rect 325660 3788 325666 3800
rect 357802 3788 357808 3800
rect 325660 3760 357808 3788
rect 325660 3748 325666 3760
rect 357802 3748 357808 3760
rect 357860 3748 357866 3800
rect 408402 3748 408408 3800
rect 408460 3788 408466 3800
rect 463970 3788 463976 3800
rect 408460 3760 463976 3788
rect 408460 3748 408466 3760
rect 463970 3748 463976 3760
rect 464028 3748 464034 3800
rect 144730 3680 144736 3732
rect 144788 3720 144794 3732
rect 179230 3720 179236 3732
rect 144788 3692 179236 3720
rect 144788 3680 144794 3692
rect 179230 3680 179236 3692
rect 179288 3680 179294 3732
rect 216582 3680 216588 3732
rect 216640 3720 216646 3732
rect 258258 3720 258264 3732
rect 216640 3692 258264 3720
rect 216640 3680 216646 3692
rect 258258 3680 258264 3692
rect 258316 3680 258322 3732
rect 322106 3680 322112 3732
rect 322164 3720 322170 3732
rect 356882 3720 356888 3732
rect 322164 3692 356888 3720
rect 322164 3680 322170 3692
rect 356882 3680 356888 3692
rect 356940 3680 356946 3732
rect 418890 3680 418896 3732
rect 418948 3720 418954 3732
rect 481726 3720 481732 3732
rect 418948 3692 481732 3720
rect 418948 3680 418954 3692
rect 481726 3680 481732 3692
rect 481784 3680 481790 3732
rect 137646 3612 137652 3664
rect 137704 3652 137710 3664
rect 182910 3652 182916 3664
rect 137704 3624 182916 3652
rect 137704 3612 137710 3624
rect 182910 3612 182916 3624
rect 182968 3612 182974 3664
rect 194410 3612 194416 3664
rect 194468 3652 194474 3664
rect 214558 3652 214564 3664
rect 194468 3624 214564 3652
rect 194468 3612 194474 3624
rect 214558 3612 214564 3624
rect 214616 3612 214622 3664
rect 216490 3612 216496 3664
rect 216548 3652 216554 3664
rect 261754 3652 261760 3664
rect 216548 3624 261760 3652
rect 216548 3612 216554 3624
rect 261754 3612 261760 3624
rect 261812 3612 261818 3664
rect 318518 3612 318524 3664
rect 318576 3652 318582 3664
rect 361666 3652 361672 3664
rect 318576 3624 361672 3652
rect 318576 3612 318582 3624
rect 361666 3612 361672 3624
rect 361724 3612 361730 3664
rect 406378 3612 406384 3664
rect 406436 3652 406442 3664
rect 478138 3652 478144 3664
rect 406436 3624 478144 3652
rect 406436 3612 406442 3624
rect 478138 3612 478144 3624
rect 478196 3612 478202 3664
rect 134150 3544 134156 3596
rect 134208 3584 134214 3596
rect 181346 3584 181352 3596
rect 134208 3556 181352 3584
rect 134208 3544 134214 3556
rect 181346 3544 181352 3556
rect 181404 3544 181410 3596
rect 190822 3544 190828 3596
rect 190880 3584 190886 3596
rect 213178 3584 213184 3596
rect 190880 3556 213184 3584
rect 190880 3544 190886 3556
rect 213178 3544 213184 3556
rect 213236 3544 213242 3596
rect 219066 3544 219072 3596
rect 219124 3584 219130 3596
rect 265342 3584 265348 3596
rect 219124 3556 265348 3584
rect 219124 3544 219130 3556
rect 265342 3544 265348 3556
rect 265400 3544 265406 3596
rect 315022 3544 315028 3596
rect 315080 3584 315086 3596
rect 358906 3584 358912 3596
rect 315080 3556 358912 3584
rect 315080 3544 315086 3556
rect 358906 3544 358912 3556
rect 358964 3544 358970 3596
rect 381538 3544 381544 3596
rect 381596 3584 381602 3596
rect 474550 3584 474556 3596
rect 381596 3556 474556 3584
rect 381596 3544 381602 3556
rect 474550 3544 474556 3556
rect 474608 3544 474614 3596
rect 565078 3544 565084 3596
rect 565136 3584 565142 3596
rect 573910 3584 573916 3596
rect 565136 3556 573916 3584
rect 565136 3544 565142 3556
rect 573910 3544 573916 3556
rect 573968 3544 573974 3596
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 205634 3516 205640 3528
rect 148376 3488 205640 3516
rect 148376 3476 148382 3488
rect 205634 3476 205640 3488
rect 205692 3476 205698 3528
rect 219986 3476 219992 3528
rect 220044 3516 220050 3528
rect 268838 3516 268844 3528
rect 220044 3488 268844 3516
rect 220044 3476 220050 3488
rect 268838 3476 268844 3488
rect 268896 3476 268902 3528
rect 311434 3476 311440 3528
rect 311492 3516 311498 3528
rect 358998 3516 359004 3528
rect 311492 3488 359004 3516
rect 311492 3476 311498 3488
rect 358998 3476 359004 3488
rect 359056 3476 359062 3528
rect 398834 3476 398840 3528
rect 398892 3516 398898 3528
rect 400122 3516 400128 3528
rect 398892 3488 400128 3516
rect 398892 3476 398898 3488
rect 400122 3476 400128 3488
rect 400180 3476 400186 3528
rect 416498 3476 416504 3528
rect 416556 3516 416562 3528
rect 417878 3516 417884 3528
rect 416556 3488 417884 3516
rect 416556 3476 416562 3488
rect 417878 3476 417884 3488
rect 417936 3476 417942 3528
rect 510062 3516 510068 3528
rect 417988 3488 510068 3516
rect 141234 3408 141240 3460
rect 141292 3448 141298 3460
rect 202874 3448 202880 3460
rect 141292 3420 202880 3448
rect 141292 3408 141298 3420
rect 202874 3408 202880 3420
rect 202932 3408 202938 3460
rect 205082 3408 205088 3460
rect 205140 3448 205146 3460
rect 215938 3448 215944 3460
rect 205140 3420 215944 3448
rect 205140 3408 205146 3420
rect 215938 3408 215944 3420
rect 215996 3408 216002 3460
rect 219894 3408 219900 3460
rect 219952 3448 219958 3460
rect 272426 3448 272432 3460
rect 219952 3420 272432 3448
rect 219952 3408 219958 3420
rect 272426 3408 272432 3420
rect 272484 3408 272490 3460
rect 307938 3408 307944 3460
rect 307996 3448 308002 3460
rect 356606 3448 356612 3460
rect 307996 3420 356612 3448
rect 307996 3408 308002 3420
rect 356606 3408 356612 3420
rect 356664 3408 356670 3460
rect 359642 3408 359648 3460
rect 359700 3448 359706 3460
rect 359700 3420 412634 3448
rect 359700 3408 359706 3420
rect 217502 3340 217508 3392
rect 217560 3380 217566 3392
rect 233418 3380 233424 3392
rect 217560 3352 233424 3380
rect 217560 3340 217566 3352
rect 233418 3340 233424 3352
rect 233476 3340 233482 3392
rect 346946 3340 346952 3392
rect 347004 3380 347010 3392
rect 359274 3380 359280 3392
rect 347004 3352 359280 3380
rect 347004 3340 347010 3352
rect 359274 3340 359280 3352
rect 359332 3340 359338 3392
rect 217594 3272 217600 3324
rect 217652 3312 217658 3324
rect 229830 3312 229836 3324
rect 217652 3284 229836 3312
rect 217652 3272 217658 3284
rect 229830 3272 229836 3284
rect 229888 3272 229894 3324
rect 350442 3272 350448 3324
rect 350500 3312 350506 3324
rect 359090 3312 359096 3324
rect 350500 3284 359096 3312
rect 350500 3272 350506 3284
rect 359090 3272 359096 3284
rect 359148 3272 359154 3324
rect 216398 3204 216404 3256
rect 216456 3244 216462 3256
rect 226334 3244 226340 3256
rect 216456 3216 226340 3244
rect 216456 3204 216462 3216
rect 226334 3204 226340 3216
rect 226392 3204 226398 3256
rect 354030 3204 354036 3256
rect 354088 3244 354094 3256
rect 358814 3244 358820 3256
rect 354088 3216 358820 3244
rect 354088 3204 354094 3216
rect 358814 3204 358820 3216
rect 358872 3204 358878 3256
rect 412606 3244 412634 3420
rect 414842 3340 414848 3392
rect 414900 3380 414906 3392
rect 417988 3380 418016 3488
rect 510062 3476 510068 3488
rect 510120 3476 510126 3528
rect 569218 3476 569224 3528
rect 569276 3516 569282 3528
rect 577406 3516 577412 3528
rect 569276 3488 577412 3516
rect 569276 3476 569282 3488
rect 577406 3476 577412 3488
rect 577464 3476 577470 3528
rect 492306 3448 492312 3460
rect 414900 3352 418016 3380
rect 418172 3420 492312 3448
rect 414900 3340 414906 3352
rect 418172 3244 418200 3420
rect 492306 3408 492312 3420
rect 492364 3408 492370 3460
rect 562410 3408 562416 3460
rect 562468 3448 562474 3460
rect 582190 3448 582196 3460
rect 562468 3420 582196 3448
rect 562468 3408 562474 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 446214 3380 446220 3392
rect 412606 3216 418200 3244
rect 418264 3352 446220 3380
rect 415946 3136 415952 3188
rect 416004 3176 416010 3188
rect 418264 3176 418292 3352
rect 446214 3340 446220 3352
rect 446272 3340 446278 3392
rect 419074 3272 419080 3324
rect 419132 3312 419138 3324
rect 439130 3312 439136 3324
rect 419132 3284 439136 3312
rect 419132 3272 419138 3284
rect 439130 3272 439136 3284
rect 439188 3272 439194 3324
rect 418522 3204 418528 3256
rect 418580 3244 418586 3256
rect 435542 3244 435548 3256
rect 418580 3216 435548 3244
rect 418580 3204 418586 3216
rect 435542 3204 435548 3216
rect 435600 3204 435606 3256
rect 416004 3148 418292 3176
rect 416004 3136 416010 3148
rect 423674 3136 423680 3188
rect 423732 3176 423738 3188
rect 424962 3176 424968 3188
rect 423732 3148 424968 3176
rect 423732 3136 423738 3148
rect 424962 3136 424968 3148
rect 425020 3136 425026 3188
rect 578878 3068 578884 3120
rect 578936 3108 578942 3120
rect 580994 3108 581000 3120
rect 578936 3080 581000 3108
rect 578936 3068 578942 3080
rect 580994 3068 581000 3080
rect 581052 3068 581058 3120
rect 373994 2728 374000 2780
rect 374052 2768 374058 2780
rect 375282 2768 375288 2780
rect 374052 2740 375288 2768
rect 374052 2728 374058 2740
rect 375282 2728 375288 2740
rect 375340 2728 375346 2780
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 154120 700612 154172 700664
rect 163504 700612 163556 700664
rect 137836 700544 137888 700596
rect 175924 700544 175976 700596
rect 391204 700544 391256 700596
rect 429844 700544 429896 700596
rect 105452 700476 105504 700528
rect 191104 700476 191156 700528
rect 410524 700476 410576 700528
rect 494796 700476 494848 700528
rect 89168 700408 89220 700460
rect 180064 700408 180116 700460
rect 202144 700408 202196 700460
rect 235172 700408 235224 700460
rect 393964 700408 394016 700460
rect 478512 700408 478564 700460
rect 24308 700340 24360 700392
rect 166264 700340 166316 700392
rect 202236 700340 202288 700392
rect 267648 700340 267700 700392
rect 392584 700340 392636 700392
rect 527180 700340 527232 700392
rect 40500 700272 40552 700324
rect 192484 700272 192536 700324
rect 202052 700272 202104 700324
rect 283840 700272 283892 700324
rect 389824 700272 389876 700324
rect 397460 700272 397512 700324
rect 400864 700272 400916 700324
rect 559656 700272 559708 700324
rect 8116 700204 8168 700256
rect 14464 700204 14516 700256
rect 407764 699660 407816 699712
rect 413652 699660 413704 699712
rect 382924 696940 382976 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 174544 683136 174596 683188
rect 385684 683136 385736 683188
rect 580172 683136 580224 683188
rect 317420 682660 317472 682712
rect 377772 682660 377824 682712
rect 199936 682592 199988 682644
rect 221740 682592 221792 682644
rect 334164 682592 334216 682644
rect 379704 682592 379756 682644
rect 196624 682524 196676 682576
rect 255228 682524 255280 682576
rect 336556 682524 336608 682576
rect 381176 682524 381228 682576
rect 196532 682456 196584 682508
rect 276756 682456 276808 682508
rect 322204 682456 322256 682508
rect 379612 682456 379664 682508
rect 195060 682388 195112 682440
rect 279148 682388 279200 682440
rect 355692 682388 355744 682440
rect 378324 682388 378376 682440
rect 196716 682320 196768 682372
rect 281540 682320 281592 682372
rect 362868 682320 362920 682372
rect 378508 682320 378560 682372
rect 199660 682252 199712 682304
rect 226524 682252 226576 682304
rect 353300 682252 353352 682304
rect 378232 682252 378284 682304
rect 199844 682184 199896 682236
rect 231308 682184 231360 682236
rect 350908 682184 350960 682236
rect 381084 682184 381136 682236
rect 201960 682116 202012 682168
rect 236092 682116 236144 682168
rect 348516 682116 348568 682168
rect 380992 682116 381044 682168
rect 199384 682048 199436 682100
rect 233700 682048 233752 682100
rect 343732 682048 343784 682100
rect 377588 682048 377640 682100
rect 195888 681980 195940 682032
rect 252836 681980 252888 682032
rect 346124 681980 346176 682032
rect 379520 681980 379572 682032
rect 199568 681912 199620 681964
rect 212172 681912 212224 681964
rect 365260 681912 365312 681964
rect 381268 681912 381320 681964
rect 199752 681844 199804 681896
rect 216956 681844 217008 681896
rect 360476 681844 360528 681896
rect 377680 681844 377732 681896
rect 198648 681776 198700 681828
rect 219348 681776 219400 681828
rect 358084 681776 358136 681828
rect 378416 681776 378468 681828
rect 200028 681708 200080 681760
rect 207388 681708 207440 681760
rect 377220 681708 377272 681760
rect 389272 681708 389324 681760
rect 195520 680892 195572 680944
rect 257620 680892 257672 680944
rect 197084 680824 197136 680876
rect 262404 680824 262456 680876
rect 197176 680756 197228 680808
rect 267188 680756 267240 680808
rect 198464 680688 198516 680740
rect 303068 680688 303120 680740
rect 194416 680620 194468 680672
rect 307852 680620 307904 680672
rect 193036 680552 193088 680604
rect 310244 680552 310296 680604
rect 193128 680484 193180 680536
rect 312636 680484 312688 680536
rect 194508 680416 194560 680468
rect 315028 680416 315080 680468
rect 195428 680348 195480 680400
rect 329380 680348 329432 680400
rect 201684 679804 201736 679856
rect 210976 679804 211028 679856
rect 202512 679736 202564 679788
rect 206008 679736 206060 679788
rect 195152 679600 195204 679652
rect 195704 679532 195756 679584
rect 195612 679464 195664 679516
rect 195796 679396 195848 679448
rect 197268 679396 197320 679448
rect 205640 679396 205692 679448
rect 205824 679396 205876 679448
rect 206008 679396 206060 679448
rect 211114 679464 211166 679516
rect 214196 679464 214248 679516
rect 259644 679532 259696 679584
rect 223764 679464 223816 679516
rect 228548 679396 228600 679448
rect 202512 679328 202564 679380
rect 198556 679260 198608 679312
rect 201776 679260 201828 679312
rect 240508 679396 240560 679448
rect 242900 679396 242952 679448
rect 201592 679192 201644 679244
rect 202328 679192 202380 679244
rect 247684 679464 247736 679516
rect 245568 679396 245620 679448
rect 201316 679124 201368 679176
rect 201408 678988 201460 679040
rect 201684 678988 201736 679040
rect 201776 678852 201828 678904
rect 250076 679396 250128 679448
rect 324872 679396 324924 679448
rect 202328 678784 202380 678836
rect 379796 678988 379848 679040
rect 201960 678308 202012 678360
rect 202420 678308 202472 678360
rect 150992 674840 151044 674892
rect 157340 674840 157392 674892
rect 551008 674840 551060 674892
rect 557540 674840 557592 674892
rect 3516 670692 3568 670744
rect 10324 670692 10376 670744
rect 565084 670692 565136 670744
rect 580172 670692 580224 670744
rect 3424 658112 3476 658164
rect 7564 658112 7616 658164
rect 569224 643084 569276 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 573364 630640 573416 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 14556 618264 14608 618316
rect 563704 616836 563756 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 11704 605820 11756 605872
rect 403624 597524 403676 597576
rect 416780 597524 416832 597576
rect 417792 591336 417844 591388
rect 419448 591336 419500 591388
rect 558184 590656 558236 590708
rect 579804 590656 579856 590708
rect 16304 589228 16356 589280
rect 19248 589228 19300 589280
rect 51080 587800 51132 587852
rect 69756 587800 69808 587852
rect 473268 587800 473320 587852
rect 476948 587800 477000 587852
rect 522396 587800 522448 587852
rect 525892 587800 525944 587852
rect 44180 587732 44232 587784
rect 62764 587732 62816 587784
rect 50068 587664 50120 587716
rect 68652 587664 68704 587716
rect 18604 587596 18656 587648
rect 53840 587596 53892 587648
rect 55680 587596 55732 587648
rect 74356 587596 74408 587648
rect 42800 587528 42852 587580
rect 61292 587528 61344 587580
rect 414664 587528 414716 587580
rect 456064 587528 456116 587580
rect 17132 587460 17184 587512
rect 60556 587460 60608 587512
rect 79140 587460 79192 587512
rect 420000 587460 420052 587512
rect 459744 587460 459796 587512
rect 48136 587392 48188 587444
rect 66260 587392 66312 587444
rect 125968 587392 126020 587444
rect 156696 587392 156748 587444
rect 18420 587324 18472 587376
rect 39580 587324 39632 587376
rect 46848 587324 46900 587376
rect 64972 587324 65024 587376
rect 111248 587324 111300 587376
rect 162124 587324 162176 587376
rect 461584 587392 461636 587444
rect 19800 587256 19852 587308
rect 42800 587256 42852 587308
rect 16120 587188 16172 587240
rect 45284 587188 45336 587240
rect 63868 587256 63920 587308
rect 103612 587256 103664 587308
rect 156604 587256 156656 587308
rect 419908 587256 419960 587308
rect 438124 587256 438176 587308
rect 53840 587188 53892 587240
rect 73252 587188 73304 587240
rect 100944 587188 100996 587240
rect 156788 587188 156840 587240
rect 419816 587188 419868 587240
rect 439596 587188 439648 587240
rect 19984 587120 20036 587172
rect 48596 587120 48648 587172
rect 67640 587120 67692 587172
rect 98552 587120 98604 587172
rect 158076 587120 158128 587172
rect 417700 587120 417752 587172
rect 441620 587120 441672 587172
rect 16396 587052 16448 587104
rect 46848 587052 46900 587104
rect 96068 587052 96120 587104
rect 159456 587052 159508 587104
rect 413928 587052 413980 587104
rect 443092 587052 443144 587104
rect 452660 587324 452712 587376
rect 454592 587324 454644 587376
rect 473360 587324 473412 587376
rect 445668 587256 445720 587308
rect 463884 587256 463936 587308
rect 15108 586984 15160 587036
rect 44180 586984 44232 587036
rect 93584 586984 93636 587036
rect 158168 586984 158220 587036
rect 413744 586984 413796 587036
rect 444196 586984 444248 587036
rect 462780 587188 462832 587240
rect 449900 587120 449952 587172
rect 450820 587120 450872 587172
rect 459744 587120 459796 587172
rect 460664 587120 460716 587172
rect 479156 587120 479208 587172
rect 448520 587052 448572 587104
rect 467564 587052 467616 587104
rect 19708 586916 19760 586968
rect 51080 586916 51132 586968
rect 88248 586916 88300 586968
rect 159364 586916 159416 586968
rect 418804 586916 418856 586968
rect 450636 586984 450688 587036
rect 15016 586848 15068 586900
rect 48136 586848 48188 586900
rect 83648 586848 83700 586900
rect 158260 586848 158312 586900
rect 413836 586848 413888 586900
rect 445668 586848 445720 586900
rect 447324 586848 447376 586900
rect 466276 586984 466328 587036
rect 450820 586916 450872 586968
rect 468668 586916 468720 586968
rect 16488 586780 16540 586832
rect 50068 586780 50120 586832
rect 51080 586780 51132 586832
rect 52368 586780 52420 586832
rect 71136 586780 71188 586832
rect 91008 586780 91060 586832
rect 166356 586780 166408 586832
rect 445760 586780 445812 586832
rect 446496 586780 446548 586832
rect 465172 586848 465224 586900
rect 451372 586780 451424 586832
rect 469772 586780 469824 586832
rect 52644 586712 52696 586764
rect 72148 586712 72200 586764
rect 73712 586712 73764 586764
rect 157984 586712 158036 586764
rect 451280 586712 451332 586764
rect 452384 586712 452436 586764
rect 471244 586712 471296 586764
rect 15844 586644 15896 586696
rect 55680 586644 55732 586696
rect 78496 586644 78548 586696
rect 163596 586644 163648 586696
rect 419724 586644 419776 586696
rect 452660 586644 452712 586696
rect 452752 586644 452804 586696
rect 453488 586644 453540 586696
rect 16212 586576 16264 586628
rect 57060 586576 57112 586628
rect 76104 586576 76156 586628
rect 162216 586576 162268 586628
rect 416044 586576 416096 586628
rect 453580 586576 453632 586628
rect 456156 586644 456208 586696
rect 473636 586644 473688 586696
rect 472164 586576 472216 586628
rect 474096 586576 474148 586628
rect 523316 586576 523368 586628
rect 19892 586508 19944 586560
rect 36636 586508 36688 586560
rect 59820 586508 59872 586560
rect 77392 586508 77444 586560
rect 81072 586508 81124 586560
rect 167644 586508 167696 586560
rect 380164 586508 380216 586560
rect 458180 586508 458232 586560
rect 458272 586508 458324 586560
rect 478052 586508 478104 586560
rect 19248 586440 19300 586492
rect 150716 586440 150768 586492
rect 157340 586440 157392 586492
rect 417792 586440 417844 586492
rect 550824 586440 550876 586492
rect 557540 586440 557592 586492
rect 417700 586372 417752 586424
rect 449900 586372 449952 586424
rect 419356 586304 419408 586356
rect 452752 586304 452804 586356
rect 417332 586236 417384 586288
rect 451280 586236 451332 586288
rect 418620 586168 418672 586220
rect 456156 586168 456208 586220
rect 415860 586100 415912 586152
rect 456800 586100 456852 586152
rect 378968 586032 379020 586084
rect 379060 586032 379112 586084
rect 462320 586032 462372 586084
rect 470600 585964 470652 586016
rect 378968 585896 379020 585948
rect 513380 585896 513432 585948
rect 385040 585828 385092 585880
rect 522396 585828 522448 585880
rect 379060 585760 379112 585812
rect 520280 585760 520332 585812
rect 108396 585080 108448 585132
rect 200856 585080 200908 585132
rect 418896 585080 418948 585132
rect 485780 585080 485832 585132
rect 105544 585012 105596 585064
rect 200948 585012 201000 585064
rect 416596 585012 416648 585064
rect 487160 585012 487212 585064
rect 68560 584944 68612 584996
rect 197820 584944 197872 584996
rect 416504 584944 416556 584996
rect 489920 584944 489972 584996
rect 65984 584876 66036 584928
rect 197912 584876 197964 584928
rect 416228 584876 416280 584928
rect 492680 584876 492732 584928
rect 63960 584808 64012 584860
rect 198188 584808 198240 584860
rect 416688 584808 416740 584860
rect 495440 584808 495492 584860
rect 17040 584740 17092 584792
rect 59820 584740 59872 584792
rect 61844 584740 61896 584792
rect 198280 584740 198332 584792
rect 416320 584740 416372 584792
rect 498200 584740 498252 584792
rect 59268 584672 59320 584724
rect 198372 584672 198424 584724
rect 416412 584672 416464 584724
rect 500960 584672 501012 584724
rect 19064 584604 19116 584656
rect 51080 584604 51132 584656
rect 56232 584604 56284 584656
rect 198004 584604 198056 584656
rect 415952 584604 416004 584656
rect 502340 584604 502392 584656
rect 14924 584536 14976 584588
rect 52644 584536 52696 584588
rect 53656 584536 53708 584588
rect 198096 584536 198148 584588
rect 416136 584536 416188 584588
rect 505100 584536 505152 584588
rect 49792 584468 49844 584520
rect 200672 584468 200724 584520
rect 380900 584468 380952 584520
rect 474096 584468 474148 584520
rect 48688 584400 48740 584452
rect 200580 584400 200632 584452
rect 379152 584400 379204 584452
rect 510620 584400 510672 584452
rect 113824 584332 113876 584384
rect 200764 584332 200816 584384
rect 419264 584332 419316 584384
rect 483020 584332 483072 584384
rect 114560 584264 114612 584316
rect 200856 584264 200908 584316
rect 419080 584264 419132 584316
rect 480260 584264 480312 584316
rect 414848 584196 414900 584248
rect 457260 584196 457312 584248
rect 419448 583516 419500 583568
rect 445760 583516 445812 583568
rect 414756 583448 414808 583500
rect 447324 583448 447376 583500
rect 415032 583380 415084 583432
rect 448520 583380 448572 583432
rect 417240 583312 417292 583364
rect 451372 583312 451424 583364
rect 458272 583312 458324 583364
rect 414940 583244 414992 583296
rect 3332 579640 3384 579692
rect 10416 579640 10468 579692
rect 571984 576852 572036 576904
rect 580172 576852 580224 576904
rect 562324 563048 562376 563100
rect 579804 563048 579856 563100
rect 3332 553528 3384 553580
rect 7656 553528 7708 553580
rect 406384 537480 406436 537532
rect 417516 537480 417568 537532
rect 566464 536800 566516 536852
rect 580172 536800 580224 536852
rect 383016 536052 383068 536104
rect 417148 536052 417200 536104
rect 415860 535508 415912 535560
rect 416780 535508 416832 535560
rect 417884 535440 417936 535492
rect 418620 535440 418672 535492
rect 414572 533672 414624 533724
rect 417516 533672 417568 533724
rect 17408 531224 17460 531276
rect 18788 531224 18840 531276
rect 411904 530612 411956 530664
rect 416872 530612 416924 530664
rect 410616 530544 410668 530596
rect 416964 530544 417016 530596
rect 417608 530544 417660 530596
rect 16764 528572 16816 528624
rect 19340 528572 19392 528624
rect 2964 527144 3016 527196
rect 11796 527144 11848 527196
rect 570604 524424 570656 524476
rect 580172 524424 580224 524476
rect 16672 523744 16724 523796
rect 18788 523744 18840 523796
rect 16856 523676 16908 523728
rect 17776 523676 17828 523728
rect 558276 510620 558328 510672
rect 580172 510620 580224 510672
rect 17316 510552 17368 510604
rect 19248 510552 19300 510604
rect 387064 509872 387116 509924
rect 416872 509872 416924 509924
rect 389916 507832 389968 507884
rect 417792 507832 417844 507884
rect 202052 501304 202104 501356
rect 3332 500964 3384 501016
rect 15752 500964 15804 501016
rect 202236 500964 202288 501016
rect 202144 500760 202196 500812
rect 201960 500692 202012 500744
rect 207572 500692 207624 500744
rect 213368 500692 213420 500744
rect 214288 500692 214340 500744
rect 215576 500692 215628 500744
rect 215668 500692 215720 500744
rect 228364 500692 228416 500744
rect 349344 500692 349396 500744
rect 175924 500624 175976 500676
rect 216956 500624 217008 500676
rect 346400 500624 346452 500676
rect 351828 500692 351880 500744
rect 416412 500896 416464 500948
rect 416320 500828 416372 500880
rect 354864 500692 354916 500744
rect 354956 500692 355008 500744
rect 364064 500692 364116 500744
rect 364156 500692 364208 500744
rect 416688 500760 416740 500812
rect 364616 500692 364668 500744
rect 416228 500692 416280 500744
rect 196532 500556 196584 500608
rect 203064 500556 203116 500608
rect 203156 500556 203208 500608
rect 238760 500556 238812 500608
rect 343640 500556 343692 500608
rect 416504 500624 416556 500676
rect 349620 500556 349672 500608
rect 416596 500556 416648 500608
rect 174544 500488 174596 500540
rect 219440 500488 219492 500540
rect 336740 500488 336792 500540
rect 418896 500488 418948 500540
rect 196716 500420 196768 500472
rect 203156 500420 203208 500472
rect 203340 500420 203392 500472
rect 242900 500420 242952 500472
rect 333980 500420 334032 500472
rect 419264 500420 419316 500472
rect 195060 500352 195112 500404
rect 241520 500352 241572 500404
rect 329840 500352 329892 500404
rect 419080 500352 419132 500404
rect 196808 500284 196860 500336
rect 244280 500284 244332 500336
rect 327080 500284 327132 500336
rect 418988 500284 419040 500336
rect 196624 500216 196676 500268
rect 254216 500216 254268 500268
rect 324596 500216 324648 500268
rect 418712 500216 418764 500268
rect 213368 500148 213420 500200
rect 215484 500148 215536 500200
rect 340880 500148 340932 500200
rect 349620 500148 349672 500200
rect 351828 500148 351880 500200
rect 357348 500148 357400 500200
rect 357440 500148 357492 500200
rect 415952 500148 416004 500200
rect 207572 500080 207624 500132
rect 215668 500080 215720 500132
rect 351920 500080 351972 500132
rect 364064 500080 364116 500132
rect 357348 500012 357400 500064
rect 364616 500012 364668 500064
rect 19708 499944 19760 499996
rect 20628 499944 20680 499996
rect 15660 499604 15712 499656
rect 17960 499604 18012 499656
rect 15568 499536 15620 499588
rect 19708 499536 19760 499588
rect 17960 499468 18012 499520
rect 18604 499468 18656 499520
rect 244924 499468 244976 499520
rect 389916 499468 389968 499520
rect 20628 499128 20680 499180
rect 51448 499128 51500 499180
rect 18604 499060 18656 499112
rect 53840 499060 53892 499112
rect 194416 499060 194468 499112
rect 249800 499060 249852 499112
rect 17132 498992 17184 499044
rect 60740 498992 60792 499044
rect 193036 498992 193088 499044
rect 251180 498992 251232 499044
rect 7564 498924 7616 498976
rect 219532 498924 219584 498976
rect 261024 498924 261076 498976
rect 381268 498924 381320 498976
rect 17040 498856 17092 498908
rect 59544 498856 59596 498908
rect 207020 498856 207072 498908
rect 558184 498856 558236 498908
rect 19248 498788 19300 498840
rect 385776 498788 385828 498840
rect 419724 498788 419776 498840
rect 454592 498788 454644 498840
rect 15016 498448 15068 498500
rect 34520 498448 34572 498500
rect 16120 498380 16172 498432
rect 44824 498380 44876 498432
rect 45376 498380 45428 498432
rect 16028 498312 16080 498364
rect 18328 498312 18380 498364
rect 58164 498312 58216 498364
rect 15844 498244 15896 498296
rect 55864 498244 55916 498296
rect 57888 498244 57940 498296
rect 14832 498176 14884 498228
rect 15016 498176 15068 498228
rect 16304 498176 16356 498228
rect 57060 498176 57112 498228
rect 389364 498176 389416 498228
rect 389916 498176 389968 498228
rect 19064 498108 19116 498160
rect 52184 498108 52236 498160
rect 59544 498108 59596 498160
rect 78128 498108 78180 498160
rect 196440 498108 196492 498160
rect 228548 498108 228600 498160
rect 302240 498108 302292 498160
rect 413284 498108 413336 498160
rect 454592 498108 454644 498160
rect 473360 498108 473412 498160
rect 16396 498040 16448 498092
rect 46848 498040 46900 498092
rect 195520 498040 195572 498092
rect 228640 498040 228692 498092
rect 259644 498040 259696 498092
rect 378508 498040 378560 498092
rect 19984 497972 20036 498024
rect 48688 497972 48740 498024
rect 49608 497972 49660 498024
rect 195244 497972 195296 498024
rect 238852 497972 238904 498024
rect 258172 497972 258224 498024
rect 377680 497972 377732 498024
rect 18420 497904 18472 497956
rect 39672 497904 39724 497956
rect 52460 497904 52512 497956
rect 53472 497904 53524 497956
rect 71964 497904 72016 497956
rect 199200 497904 199252 497956
rect 259460 497904 259512 497956
rect 259552 497904 259604 497956
rect 379796 497904 379848 497956
rect 34520 497836 34572 497888
rect 47584 497836 47636 497888
rect 48228 497836 48280 497888
rect 51448 497836 51500 497888
rect 69664 497836 69716 497888
rect 197084 497836 197136 497888
rect 256700 497836 256752 497888
rect 258264 497836 258316 497888
rect 379612 497836 379664 497888
rect 19892 497768 19944 497820
rect 37188 497768 37240 497820
rect 42800 497768 42852 497820
rect 57888 497768 57940 497820
rect 73988 497768 74040 497820
rect 195152 497768 195204 497820
rect 255412 497768 255464 497820
rect 256792 497768 256844 497820
rect 378416 497768 378468 497820
rect 19156 497700 19208 497752
rect 36176 497700 36228 497752
rect 38660 497700 38712 497752
rect 53840 497700 53892 497752
rect 73160 497700 73212 497752
rect 201224 497700 201276 497752
rect 247132 497700 247184 497752
rect 255596 497700 255648 497752
rect 378324 497700 378376 497752
rect 445300 497700 445352 497752
rect 463700 497700 463752 497752
rect 60648 497632 60700 497684
rect 79416 497632 79468 497684
rect 196992 497632 197044 497684
rect 244372 497632 244424 497684
rect 254032 497632 254084 497684
rect 378232 497632 378284 497684
rect 419908 497632 419960 497684
rect 437480 497632 437532 497684
rect 444196 497632 444248 497684
rect 462320 497632 462372 497684
rect 462504 497632 462556 497684
rect 476120 497632 476172 497684
rect 16028 497564 16080 497616
rect 19984 497564 20036 497616
rect 22100 497564 22152 497616
rect 40592 497564 40644 497616
rect 44824 497564 44876 497616
rect 64144 497564 64196 497616
rect 196900 497564 196952 497616
rect 241612 497564 241664 497616
rect 242992 497564 243044 497616
rect 381176 497564 381228 497616
rect 419816 497564 419868 497616
rect 438860 497564 438912 497616
rect 462044 497564 462096 497616
rect 474740 497564 474792 497616
rect 19800 497496 19852 497548
rect 43444 497496 43496 497548
rect 49608 497496 49660 497548
rect 67640 497496 67692 497548
rect 68928 497496 68980 497548
rect 195336 497496 195388 497548
rect 240140 497496 240192 497548
rect 240232 497496 240284 497548
rect 379704 497496 379756 497548
rect 417976 497496 418028 497548
rect 451280 497496 451332 497548
rect 469220 497496 469272 497548
rect 15016 497428 15068 497480
rect 52460 497428 52512 497480
rect 70400 497428 70452 497480
rect 71228 497428 71280 497480
rect 313280 497428 313332 497480
rect 334900 497428 334952 497480
rect 391940 497428 391992 497480
rect 418068 497428 418120 497480
rect 452384 497428 452436 497480
rect 470876 497428 470928 497480
rect 197176 497360 197228 497412
rect 228732 497360 228784 497412
rect 360476 497360 360528 497412
rect 416136 497360 416188 497412
rect 449164 497360 449216 497412
rect 466460 497360 466512 497412
rect 450544 497292 450596 497344
rect 467840 497292 467892 497344
rect 447784 497224 447836 497276
rect 465080 497224 465132 497276
rect 20628 497156 20680 497208
rect 44180 497156 44232 497208
rect 62764 497156 62816 497208
rect 443644 497156 443696 497208
rect 461124 497156 461176 497208
rect 43444 497088 43496 497140
rect 61844 497088 61896 497140
rect 78128 497088 78180 497140
rect 79324 497088 79376 497140
rect 456064 497088 456116 497140
rect 473360 497088 473412 497140
rect 50252 497020 50304 497072
rect 68284 497020 68336 497072
rect 71964 497020 72016 497072
rect 319444 497020 319496 497072
rect 446680 497020 446732 497072
rect 465080 497020 465132 497072
rect 16488 496748 16540 496800
rect 34520 496748 34572 496800
rect 52184 496952 52236 497004
rect 52460 496952 52512 497004
rect 70400 496952 70452 497004
rect 313280 496952 313332 497004
rect 315304 496952 315356 497004
rect 459560 496952 459612 497004
rect 460572 496952 460624 497004
rect 478880 496952 478932 497004
rect 39672 496884 39724 496936
rect 44180 496884 44232 496936
rect 48228 496884 48280 496936
rect 66260 496884 66312 496936
rect 66904 496884 66956 496936
rect 68928 496884 68980 496936
rect 301504 496884 301556 496936
rect 311164 496884 311216 496936
rect 40592 496816 40644 496868
rect 43444 496816 43496 496868
rect 46848 496816 46900 496868
rect 65524 496816 65576 496868
rect 417332 496884 417384 496936
rect 418068 496884 418120 496936
rect 453304 496884 453356 496936
rect 471980 496884 472032 496936
rect 417240 496816 417292 496868
rect 417976 496816 418028 496868
rect 420736 496816 420788 496868
rect 436100 496816 436152 496868
rect 458824 496816 458876 496868
rect 459468 496816 459520 496868
rect 477500 496816 477552 496868
rect 420000 496748 420052 496800
rect 459560 496748 459612 496800
rect 15108 496680 15160 496732
rect 19800 496680 19852 496732
rect 20628 496680 20680 496732
rect 419448 496680 419500 496732
rect 445760 496680 445812 496732
rect 446680 496680 446732 496732
rect 201592 496204 201644 496256
rect 235264 496204 235316 496256
rect 212724 496136 212776 496188
rect 389824 496136 389876 496188
rect 63684 496068 63736 496120
rect 305000 496068 305052 496120
rect 316040 496068 316092 496120
rect 470784 496068 470836 496120
rect 338764 495524 338816 495576
rect 418160 495524 418212 495576
rect 420000 495524 420052 495576
rect 278044 495456 278096 495508
rect 418712 495456 418764 495508
rect 286324 495184 286376 495236
rect 413744 495184 413796 495236
rect 415308 495184 415360 495236
rect 252836 495116 252888 495168
rect 381084 495116 381136 495168
rect 248420 495048 248472 495100
rect 377588 495048 377640 495100
rect 194508 494980 194560 495032
rect 232504 494980 232556 495032
rect 249892 494980 249944 495032
rect 379520 494980 379572 495032
rect 193128 494912 193180 494964
rect 232596 494912 232648 494964
rect 251272 494912 251324 494964
rect 380992 494912 381044 494964
rect 106096 494844 106148 494896
rect 360292 494844 360344 494896
rect 415308 494844 415360 494896
rect 444196 494844 444248 494896
rect 16948 494776 17000 494828
rect 304356 494776 304408 494828
rect 319076 494776 319128 494828
rect 473544 494776 473596 494828
rect 207112 494708 207164 494760
rect 571984 494708 572036 494760
rect 48320 493484 48372 493536
rect 280252 493484 280304 493536
rect 41880 493416 41932 493468
rect 293960 493416 294012 493468
rect 325976 493416 326028 493468
rect 477592 493416 477644 493468
rect 100944 493348 100996 493400
rect 354772 493348 354824 493400
rect 208400 493280 208452 493332
rect 569224 493280 569276 493332
rect 293960 492668 294012 492720
rect 294236 492668 294288 492720
rect 416688 492668 416740 492720
rect 416780 492600 416832 492652
rect 417792 492600 417844 492652
rect 456892 492600 456944 492652
rect 208492 492056 208544 492108
rect 382924 492056 382976 492108
rect 73712 491988 73764 492040
rect 320272 491988 320324 492040
rect 328460 491988 328512 492040
rect 480536 491988 480588 492040
rect 108856 491920 108908 491972
rect 363236 491920 363288 491972
rect 329104 491308 329156 491360
rect 417792 491308 417844 491360
rect 292488 490832 292540 490884
rect 413836 490832 413888 490884
rect 415216 490832 415268 490884
rect 209780 490764 209832 490816
rect 385684 490764 385736 490816
rect 61844 490696 61896 490748
rect 281816 490696 281868 490748
rect 301044 490696 301096 490748
rect 460940 490696 460992 490748
rect 68560 490628 68612 490680
rect 313280 490628 313332 490680
rect 415216 490628 415268 490680
rect 445300 490628 445352 490680
rect 76840 490560 76892 490612
rect 322940 490560 322992 490612
rect 342260 490560 342312 490612
rect 490472 490560 490524 490612
rect 64144 489812 64196 489864
rect 291200 489812 291252 489864
rect 159456 489268 159508 489320
rect 349252 489268 349304 489320
rect 37280 489200 37332 489252
rect 280804 489200 280856 489252
rect 287060 489200 287112 489252
rect 452660 489200 452712 489252
rect 78588 489132 78640 489184
rect 325792 489132 325844 489184
rect 353300 489132 353352 489184
rect 500960 489132 501012 489184
rect 291200 488724 291252 488776
rect 292488 488724 292540 488776
rect 417884 488452 417936 488504
rect 456064 488452 456116 488504
rect 292856 487976 292908 488028
rect 455512 487976 455564 488028
rect 158260 487908 158312 487960
rect 334072 487908 334124 487960
rect 66904 487840 66956 487892
rect 300124 487840 300176 487892
rect 88248 487772 88300 487824
rect 339500 487772 339552 487824
rect 350540 487772 350592 487824
rect 497464 487772 497516 487824
rect 324504 487160 324556 487212
rect 415124 487160 415176 487212
rect 417884 487160 417936 487212
rect 62764 487092 62816 487144
rect 286324 487092 286376 487144
rect 282920 486616 282972 486668
rect 449900 486616 449952 486668
rect 158168 486548 158220 486600
rect 346492 486548 346544 486600
rect 91008 486480 91060 486532
rect 342352 486480 342404 486532
rect 208584 486412 208636 486464
rect 573364 486412 573416 486464
rect 285680 485868 285732 485920
rect 286324 485868 286376 485920
rect 73988 485732 74040 485784
rect 324504 485732 324556 485784
rect 156788 485188 156840 485240
rect 356060 485188 356112 485240
rect 10324 485120 10376 485172
rect 221096 485120 221148 485172
rect 96528 485052 96580 485104
rect 347780 485052 347832 485104
rect 209044 484372 209096 484424
rect 580172 484372 580224 484424
rect 281816 484304 281868 484356
rect 413928 484304 413980 484356
rect 417884 484304 417936 484356
rect 163596 483828 163648 483880
rect 327172 483828 327224 483880
rect 417884 483828 417936 483880
rect 443644 483828 443696 483880
rect 3424 483760 3476 483812
rect 222476 483760 222528 483812
rect 296904 483760 296956 483812
rect 458180 483760 458232 483812
rect 86868 483692 86920 483744
rect 336832 483692 336884 483744
rect 345020 483692 345072 483744
rect 492680 483692 492732 483744
rect 205640 483624 205692 483676
rect 570604 483624 570656 483676
rect 305092 482468 305144 482520
rect 462412 482468 462464 482520
rect 71688 482400 71740 482452
rect 316132 482400 316184 482452
rect 84108 482332 84160 482384
rect 332600 482332 332652 482384
rect 338120 482332 338172 482384
rect 487160 482332 487212 482384
rect 205732 482264 205784 482316
rect 566464 482264 566516 482316
rect 415032 481584 415084 481636
rect 449164 481584 449216 481636
rect 201500 481040 201552 481092
rect 215576 481040 215628 481092
rect 309140 481040 309192 481092
rect 465172 481040 465224 481092
rect 66168 480972 66220 481024
rect 309232 480972 309284 481024
rect 81348 480904 81400 480956
rect 329932 480904 329984 480956
rect 335360 480904 335412 480956
rect 485780 480904 485832 480956
rect 301504 480224 301556 480276
rect 415032 480224 415084 480276
rect 319444 480156 319496 480208
rect 419356 480156 419408 480208
rect 278780 479612 278832 479664
rect 447140 479612 447192 479664
rect 159364 479544 159416 479596
rect 340972 479544 341024 479596
rect 93768 479476 93820 479528
rect 345112 479476 345164 479528
rect 419356 479476 419408 479528
rect 420000 479476 420052 479528
rect 453304 479476 453356 479528
rect 318892 478864 318944 478916
rect 319444 478864 319496 478916
rect 104808 478252 104860 478304
rect 357532 478252 357584 478304
rect 19432 478184 19484 478236
rect 295340 478184 295392 478236
rect 332692 478184 332744 478236
rect 483020 478184 483072 478236
rect 205824 478116 205876 478168
rect 562324 478116 562376 478168
rect 68284 476892 68336 476944
rect 307024 476892 307076 476944
rect 115848 476824 115900 476876
rect 371240 476824 371292 476876
rect 19340 476756 19392 476808
rect 311900 476756 311952 476808
rect 321560 476756 321612 476808
rect 476120 476756 476172 476808
rect 209964 475532 210016 475584
rect 392584 475532 392636 475584
rect 11704 475464 11756 475516
rect 220912 475464 220964 475516
rect 287152 475464 287204 475516
rect 403624 475464 403676 475516
rect 73804 475396 73856 475448
rect 322204 475396 322256 475448
rect 99288 475328 99340 475380
rect 352012 475328 352064 475380
rect 356152 475328 356204 475380
rect 502340 475328 502392 475380
rect 3056 474716 3108 474768
rect 80704 474716 80756 474768
rect 303804 474172 303856 474224
rect 417424 474172 417476 474224
rect 43444 474104 43496 474156
rect 290464 474104 290516 474156
rect 294052 474104 294104 474156
rect 414664 474104 414716 474156
rect 114468 474036 114520 474088
rect 368756 474036 368808 474088
rect 379520 474036 379572 474088
rect 523040 474036 523092 474088
rect 205916 473968 205968 474020
rect 558276 473968 558328 474020
rect 405648 473288 405700 473340
rect 406384 473288 406436 473340
rect 162216 472812 162268 472864
rect 324504 472812 324556 472864
rect 158076 472744 158128 472796
rect 353392 472744 353444 472796
rect 76564 472676 76616 472728
rect 331220 472676 331272 472728
rect 17684 472608 17736 472660
rect 308496 472608 308548 472660
rect 358820 472608 358872 472660
rect 504364 472608 504416 472660
rect 311900 471996 311952 472048
rect 405648 471996 405700 472048
rect 75184 471928 75236 471980
rect 328552 471928 328604 471980
rect 329104 471928 329156 471980
rect 414848 471928 414900 471980
rect 457444 471928 457496 471980
rect 166264 471384 166316 471436
rect 219624 471384 219676 471436
rect 331220 471384 331272 471436
rect 414848 471384 414900 471436
rect 166356 471316 166408 471368
rect 343732 471316 343784 471368
rect 53748 471248 53800 471300
rect 288532 471248 288584 471300
rect 311992 471248 312044 471300
rect 467932 471248 467984 471300
rect 204260 470568 204312 470620
rect 579988 470568 580040 470620
rect 69664 470500 69716 470552
rect 311164 470500 311216 470552
rect 417700 470500 417752 470552
rect 450544 470500 450596 470552
rect 118608 469888 118660 469940
rect 375380 469888 375432 469940
rect 17592 469820 17644 469872
rect 300768 469820 300820 469872
rect 371332 469820 371384 469872
rect 514760 469820 514812 469872
rect 307024 469344 307076 469396
rect 310520 469276 310572 469328
rect 311164 469276 311216 469328
rect 417700 469276 417752 469328
rect 303712 469208 303764 469260
rect 304356 469208 304408 469260
rect 413928 469208 413980 469260
rect 414572 469208 414624 469260
rect 300768 469140 300820 469192
rect 407856 469140 407908 469192
rect 414756 469140 414808 469192
rect 447784 469140 447836 469192
rect 201316 468664 201368 468716
rect 252652 468664 252704 468716
rect 300124 468664 300176 468716
rect 414572 468664 414624 468716
rect 414756 468664 414808 468716
rect 197268 468596 197320 468648
rect 249984 468596 250036 468648
rect 284484 468596 284536 468648
rect 418804 468596 418856 468648
rect 167644 468528 167696 468580
rect 331312 468528 331364 468580
rect 16856 468460 16908 468512
rect 295432 468460 295484 468512
rect 363052 468460 363104 468512
rect 507860 468460 507912 468512
rect 299480 467848 299532 467900
rect 300124 467848 300176 467900
rect 313372 467236 313424 467288
rect 388444 467236 388496 467288
rect 157984 467168 158036 467220
rect 321652 467168 321704 467220
rect 16672 467100 16724 467152
rect 291292 467100 291344 467152
rect 368572 467100 368624 467152
rect 512644 467100 512696 467152
rect 295432 466488 295484 466540
rect 19064 466420 19116 466472
rect 42800 466420 42852 466472
rect 43628 466420 43680 466472
rect 79416 466420 79468 466472
rect 80060 466420 80112 466472
rect 338304 466420 338356 466472
rect 338764 466420 338816 466472
rect 411168 466420 411220 466472
rect 411904 466420 411956 466472
rect 198648 466352 198700 466404
rect 241704 466352 241756 466404
rect 411260 466352 411312 466404
rect 414940 466352 414992 466404
rect 458824 466352 458876 466404
rect 202420 466284 202472 466336
rect 248512 466284 248564 466336
rect 195704 466216 195756 466268
rect 243084 466216 243136 466268
rect 199384 466148 199436 466200
rect 247224 466148 247276 466200
rect 195612 466080 195664 466132
rect 245844 466080 245896 466132
rect 202328 466012 202380 466064
rect 252744 466012 252796 466064
rect 198556 465944 198608 465996
rect 251364 465944 251416 465996
rect 195796 465876 195848 465928
rect 250076 465876 250128 465928
rect 197912 465808 197964 465860
rect 310612 465808 310664 465860
rect 43628 465740 43680 465792
rect 281724 465740 281776 465792
rect 301504 465740 301556 465792
rect 304264 465740 304316 465792
rect 365904 465740 365956 465792
rect 510620 465740 510672 465792
rect 126888 465672 126940 465724
rect 383660 465672 383712 465724
rect 201408 465604 201460 465656
rect 240324 465604 240376 465656
rect 65524 465536 65576 465588
rect 66260 465536 66312 465588
rect 199292 465536 199344 465588
rect 237472 465536 237524 465588
rect 409788 465536 409840 465588
rect 410616 465536 410668 465588
rect 291292 465128 291344 465180
rect 409788 465128 409840 465180
rect 18972 465060 19024 465112
rect 38660 465060 38712 465112
rect 66260 465060 66312 465112
rect 295708 465060 295760 465112
rect 336648 465060 336700 465112
rect 411260 465060 411312 465112
rect 412548 465060 412600 465112
rect 277492 464992 277544 465044
rect 278044 464992 278096 465044
rect 287704 464992 287756 465044
rect 288348 464992 288400 465044
rect 415860 464992 415912 465044
rect 417424 464992 417476 465044
rect 440240 464992 440292 465044
rect 79324 464924 79376 464976
rect 80152 464924 80204 464976
rect 187608 464448 187660 464500
rect 232688 464448 232740 464500
rect 290464 464448 290516 464500
rect 417424 464448 417476 464500
rect 186872 464380 186924 464432
rect 232780 464380 232832 464432
rect 374000 464380 374052 464432
rect 517520 464380 517572 464432
rect 124128 464312 124180 464364
rect 380992 464312 381044 464364
rect 188988 464244 189040 464296
rect 235356 464244 235408 464296
rect 191472 464176 191524 464228
rect 273352 464176 273404 464228
rect 289820 464176 289872 464228
rect 290464 464176 290516 464228
rect 188160 464108 188212 464160
rect 271880 464108 271932 464160
rect 186780 464040 186832 464092
rect 271972 464040 272024 464092
rect 183468 463972 183520 464024
rect 270776 463972 270828 464024
rect 186228 463904 186280 463956
rect 274732 463904 274784 463956
rect 184848 463836 184900 463888
rect 274824 463836 274876 463888
rect 186136 463768 186188 463820
rect 276204 463768 276256 463820
rect 18880 463700 18932 463752
rect 44180 463700 44232 463752
rect 44640 463700 44692 463752
rect 80152 463700 80204 463752
rect 335452 463700 335504 463752
rect 336648 463700 336700 463752
rect 199752 463632 199804 463684
rect 241796 463632 241848 463684
rect 308496 463632 308548 463684
rect 309048 463632 309100 463684
rect 383016 463632 383068 463684
rect 199936 463564 199988 463616
rect 243176 463564 243228 463616
rect 199660 463496 199712 463548
rect 244556 463496 244608 463548
rect 199844 463428 199896 463480
rect 247316 463428 247368 463480
rect 195888 463360 195940 463412
rect 254124 463360 254176 463412
rect 200580 463292 200632 463344
rect 281632 463292 281684 463344
rect 200672 463224 200724 463276
rect 285772 463224 285824 463276
rect 200948 463156 201000 463208
rect 361580 463156 361632 463208
rect 201040 463088 201092 463140
rect 364340 463088 364392 463140
rect 419448 463088 419500 463140
rect 436192 463088 436244 463140
rect 44640 463020 44692 463072
rect 285864 463020 285916 463072
rect 376760 463020 376812 463072
rect 519544 463020 519596 463072
rect 121368 462952 121420 463004
rect 378232 462952 378284 463004
rect 414756 462952 414808 463004
rect 445760 462952 445812 463004
rect 199568 462884 199620 462936
rect 239036 462884 239088 462936
rect 199476 462816 199528 462868
rect 236184 462816 236236 462868
rect 295708 462408 295760 462460
rect 414756 462408 414808 462460
rect 3424 462340 3476 462392
rect 218060 462340 218112 462392
rect 281724 462340 281776 462392
rect 419448 462340 419500 462392
rect 192484 461932 192536 461984
rect 218152 461932 218204 461984
rect 191104 461864 191156 461916
rect 216772 461864 216824 461916
rect 169760 461796 169812 461848
rect 216864 461796 216916 461848
rect 218060 461796 218112 461848
rect 225052 461796 225104 461848
rect 200856 461728 200908 461780
rect 374092 461728 374144 461780
rect 14464 461660 14516 461712
rect 219716 461660 219768 461712
rect 298284 461660 298336 461712
rect 380164 461660 380216 461712
rect 10416 461592 10468 461644
rect 222292 461592 222344 461644
rect 347872 461592 347924 461644
rect 494704 461592 494756 461644
rect 191748 461388 191800 461440
rect 270592 461388 270644 461440
rect 185860 461320 185912 461372
rect 266360 461320 266412 461372
rect 189540 461252 189592 461304
rect 270684 461252 270736 461304
rect 190368 461184 190420 461236
rect 272064 461184 272116 461236
rect 185768 461116 185820 461168
rect 267740 461116 267792 461168
rect 173624 461048 173676 461100
rect 294144 461048 294196 461100
rect 173440 460980 173492 461032
rect 306380 460980 306432 461032
rect 198740 460912 198792 460964
rect 580632 460912 580684 460964
rect 385776 460844 385828 460896
rect 387064 460844 387116 460896
rect 200028 460640 200080 460692
rect 237932 460640 237984 460692
rect 198096 460572 198148 460624
rect 290188 460572 290240 460624
rect 198004 460504 198056 460556
rect 294604 460504 294656 460556
rect 198372 460436 198424 460488
rect 299020 460436 299072 460488
rect 198280 460368 198332 460420
rect 303068 460368 303120 460420
rect 198188 460300 198240 460352
rect 307116 460300 307168 460352
rect 156604 460232 156656 460284
rect 358912 460232 358964 460284
rect 3608 460164 3660 460216
rect 223948 460164 224000 460216
rect 185952 459892 186004 459944
rect 269120 459892 269172 459944
rect 186044 459824 186096 459876
rect 276112 459824 276164 459876
rect 181444 459756 181496 459808
rect 280988 459756 281040 459808
rect 181720 459688 181772 459740
rect 301228 459688 301280 459740
rect 179052 459620 179104 459672
rect 324320 459620 324372 459672
rect 181628 459552 181680 459604
rect 381084 459552 381136 459604
rect 374000 459484 374052 459536
rect 374460 459484 374512 459536
rect 181536 459212 181588 459264
rect 321100 459212 321152 459264
rect 178776 459144 178828 459196
rect 327724 459144 327776 459196
rect 180064 459076 180116 459128
rect 218428 459076 218480 459128
rect 163504 459008 163556 459060
rect 216680 459008 216732 459060
rect 188620 458940 188672 458992
rect 262956 458940 263008 458992
rect 15752 458872 15804 458924
rect 223672 458872 223724 458924
rect 7656 458804 7708 458856
rect 222476 458804 222528 458856
rect 190276 458736 190328 458788
rect 267004 458736 267056 458788
rect 306012 458736 306064 458788
rect 402244 458736 402296 458788
rect 184756 458668 184808 458720
rect 277584 458668 277636 458720
rect 302516 458668 302568 458720
rect 402336 458668 402388 458720
rect 310060 458600 310112 458652
rect 399668 458600 399720 458652
rect 313740 458532 313792 458584
rect 399484 458532 399536 458584
rect 181904 458464 181956 458516
rect 313188 458464 313240 458516
rect 317052 458464 317104 458516
rect 399576 458464 399628 458516
rect 178684 458396 178736 458448
rect 334348 458396 334400 458448
rect 178868 458328 178920 458380
rect 341064 458328 341116 458380
rect 198832 458260 198884 458312
rect 580448 458260 580500 458312
rect 199292 458192 199344 458244
rect 580724 458192 580776 458244
rect 80704 457784 80756 457836
rect 224316 457784 224368 457836
rect 353300 457784 353352 457836
rect 353852 457784 353904 457836
rect 210056 457716 210108 457768
rect 400864 457716 400916 457768
rect 14556 457648 14608 457700
rect 221004 457648 221056 457700
rect 4804 457580 4856 457632
rect 220820 457580 220872 457632
rect 208860 457512 208912 457564
rect 565084 457512 565136 457564
rect 207756 457444 207808 457496
rect 563704 457444 563756 457496
rect 201500 457308 201552 457360
rect 209136 457308 209188 457360
rect 191656 457240 191708 457292
rect 264980 457240 265032 457292
rect 186964 457172 187016 457224
rect 319628 457172 319680 457224
rect 187056 457104 187108 457156
rect 326252 457104 326304 457156
rect 184204 457036 184256 457088
rect 360200 457036 360252 457088
rect 184296 456968 184348 457020
rect 365996 456968 366048 457020
rect 204352 456900 204404 456952
rect 394148 456900 394200 456952
rect 203064 456832 203116 456884
rect 399760 456832 399812 456884
rect 204812 456764 204864 456816
rect 209044 456764 209096 456816
rect 209136 456764 209188 456816
rect 403624 456764 403676 456816
rect 200672 456424 200724 456476
rect 209504 456424 209556 456476
rect 181996 456356 182048 456408
rect 293040 456356 293092 456408
rect 183376 456288 183428 456340
rect 269948 456288 270000 456340
rect 310520 456288 310572 456340
rect 311532 456288 311584 456340
rect 322204 456288 322256 456340
rect 419632 456288 419684 456340
rect 187240 456220 187292 456272
rect 279516 456220 279568 456272
rect 285864 456220 285916 456272
rect 286140 456220 286192 456272
rect 286600 456220 286652 456272
rect 287060 456220 287112 456272
rect 287980 456220 288032 456272
rect 288440 456220 288492 456272
rect 289452 456220 289504 456272
rect 303620 456220 303672 456272
rect 304264 456220 304316 456272
rect 305000 456220 305052 456272
rect 305644 456220 305696 456272
rect 310612 456220 310664 456272
rect 311164 456220 311216 456272
rect 317328 456220 317380 456272
rect 323216 456220 323268 456272
rect 419540 456220 419592 456272
rect 437480 456220 437532 456272
rect 162124 456152 162176 456204
rect 367836 456152 367888 456204
rect 379520 456152 379572 456204
rect 380348 456152 380400 456204
rect 380900 456152 380952 456204
rect 381820 456152 381872 456204
rect 386144 456152 386196 456204
rect 387064 456152 387116 456204
rect 11796 456084 11848 456136
rect 222200 456084 222252 456136
rect 254032 456084 254084 456136
rect 254492 456084 254544 456136
rect 255412 456084 255464 456136
rect 256332 456084 256384 456136
rect 258172 456084 258224 456136
rect 258540 456084 258592 456136
rect 270684 456084 270736 456136
rect 271420 456084 271472 456136
rect 271880 456084 271932 456136
rect 272524 456084 272576 456136
rect 273260 456084 273312 456136
rect 273996 456084 274048 456136
rect 277400 456084 277452 456136
rect 278412 456084 278464 456136
rect 280160 456084 280212 456136
rect 280620 456084 280672 456136
rect 281724 456084 281776 456136
rect 282460 456084 282512 456136
rect 285680 456084 285732 456136
rect 286508 456084 286560 456136
rect 286600 456084 286652 456136
rect 419724 456152 419776 456204
rect 438860 456152 438912 456204
rect 419632 456084 419684 456136
rect 419908 456084 419960 456136
rect 454684 456084 454736 456136
rect 205640 456016 205692 456068
rect 206284 456016 206336 456068
rect 208492 456016 208544 456068
rect 209228 456016 209280 456068
rect 209320 456016 209372 456068
rect 580172 456016 580224 456068
rect 187148 455948 187200 456000
rect 317328 455948 317380 456000
rect 317420 455948 317472 456000
rect 318156 455948 318208 456000
rect 320180 455948 320232 456000
rect 320732 455948 320784 456000
rect 331220 455948 331272 456000
rect 331772 455948 331824 456000
rect 332600 455948 332652 456000
rect 333244 455948 333296 456000
rect 335360 455948 335412 456000
rect 335820 455948 335872 456000
rect 336740 455948 336792 456000
rect 337292 455948 337344 456000
rect 338120 455948 338172 456000
rect 339132 455948 339184 456000
rect 347780 455948 347832 456000
rect 348700 455948 348752 456000
rect 351920 455948 351972 456000
rect 352380 455948 352432 456000
rect 354680 455948 354732 456000
rect 355324 455948 355376 456000
rect 357440 455948 357492 456000
rect 358268 455948 358320 456000
rect 364340 455948 364392 456000
rect 364892 455948 364944 456000
rect 205824 455880 205876 455932
rect 206652 455880 206704 455932
rect 209872 455880 209924 455932
rect 210700 455880 210752 455932
rect 211252 455880 211304 455932
rect 212172 455880 212224 455932
rect 280804 455880 280856 455932
rect 419540 455880 419592 455932
rect 419816 455880 419868 455932
rect 184480 455812 184532 455864
rect 363144 455812 363196 455864
rect 184388 455744 184440 455796
rect 368940 455744 368992 455796
rect 204720 455676 204772 455728
rect 209320 455676 209372 455728
rect 209412 455676 209464 455728
rect 391296 455676 391348 455728
rect 202512 455608 202564 455660
rect 395436 455608 395488 455660
rect 201776 455540 201828 455592
rect 209412 455540 209464 455592
rect 209504 455540 209556 455592
rect 395344 455540 395396 455592
rect 201040 455472 201092 455524
rect 396724 455472 396776 455524
rect 198464 455404 198516 455456
rect 562324 455404 562376 455456
rect 157984 454996 158036 455048
rect 367468 454996 367520 455048
rect 181352 454928 181404 454980
rect 227996 454928 228048 454980
rect 184020 454860 184072 454912
rect 227260 454860 227312 454912
rect 368756 454860 368808 454912
rect 402520 454860 402572 454912
rect 188712 454792 188764 454844
rect 262588 454792 262640 454844
rect 357900 454792 357952 454844
rect 402796 454792 402848 454844
rect 188804 454724 188856 454776
rect 264060 454724 264112 454776
rect 343180 454724 343232 454776
rect 405096 454724 405148 454776
rect 111708 454656 111760 454708
rect 366364 454656 366416 454708
rect 383292 454656 383344 454708
rect 525800 454656 525852 454708
rect 187516 454588 187568 454640
rect 268108 454588 268160 454640
rect 333612 454588 333664 454640
rect 405004 454588 405056 454640
rect 202880 454520 202932 454572
rect 390284 454520 390336 454572
rect 200304 454452 200356 454504
rect 392676 454452 392728 454504
rect 199200 454384 199252 454436
rect 394056 454384 394108 454436
rect 354956 454316 355008 454368
rect 402704 454316 402756 454368
rect 14464 454248 14516 454300
rect 233884 454248 233936 454300
rect 327264 454248 327316 454300
rect 407764 454248 407816 454300
rect 10324 454180 10376 454232
rect 231308 454180 231360 454232
rect 323952 454180 324004 454232
rect 407948 454180 408000 454232
rect 7564 454112 7616 454164
rect 233516 454112 233568 454164
rect 293776 454112 293828 454164
rect 410524 454112 410576 454164
rect 198096 454044 198148 454096
rect 570604 454044 570656 454096
rect 280528 453636 280580 453688
rect 393964 453636 394016 453688
rect 200856 453568 200908 453620
rect 371056 453568 371108 453620
rect 50988 453500 51040 453552
rect 284576 453500 284628 453552
rect 56508 453432 56560 453484
rect 293408 453432 293460 453484
rect 361120 453432 361172 453484
rect 402612 453432 402664 453484
rect 59268 453364 59320 453416
rect 297824 453364 297876 453416
rect 362592 453364 362644 453416
rect 410708 453364 410760 453416
rect 62028 453296 62080 453348
rect 301872 453296 301924 453348
rect 346400 453296 346452 453348
rect 405280 453296 405332 453348
rect 337200 453228 337252 453280
rect 405372 453228 405424 453280
rect 193864 453160 193916 453212
rect 224960 453160 225012 453212
rect 324320 453160 324372 453212
rect 324688 453160 324740 453212
rect 344928 453160 344980 453212
rect 413376 453160 413428 453212
rect 191012 453092 191064 453144
rect 229744 453092 229796 453144
rect 240232 453092 240284 453144
rect 240876 453092 240928 453144
rect 241612 453092 241664 453144
rect 242348 453092 242400 453144
rect 245752 453092 245804 453144
rect 246396 453092 246448 453144
rect 247040 453092 247092 453144
rect 247868 453092 247920 453144
rect 324504 453092 324556 453144
rect 324780 453092 324832 453144
rect 330576 453092 330628 453144
rect 405188 453092 405240 453144
rect 185400 453024 185452 453076
rect 229376 453024 229428 453076
rect 237472 453024 237524 453076
rect 238300 453024 238352 453076
rect 238760 453024 238812 453076
rect 239404 453024 239456 453076
rect 240140 453024 240192 453076
rect 240600 453024 240652 453076
rect 241704 453024 241756 453076
rect 241980 453024 242032 453076
rect 243084 453024 243136 453076
rect 243820 453024 243872 453076
rect 244280 453024 244332 453076
rect 244924 453024 244976 453076
rect 245660 453024 245712 453076
rect 246120 453024 246172 453076
rect 247224 453024 247276 453076
rect 247500 453024 247552 453076
rect 249984 453024 250036 453076
rect 250812 453024 250864 453076
rect 252744 453024 252796 453076
rect 253388 453024 253440 453076
rect 295432 453024 295484 453076
rect 295800 453024 295852 453076
rect 315856 453024 315908 453076
rect 407856 453024 407908 453076
rect 188436 452956 188488 453008
rect 262128 452956 262180 453008
rect 295340 452956 295392 453008
rect 296076 452956 296128 453008
rect 321560 452956 321612 453008
rect 322572 452956 322624 453008
rect 324412 452956 324464 453008
rect 325148 452956 325200 453008
rect 325792 452956 325844 453008
rect 326620 452956 326672 453008
rect 328460 452956 328512 453008
rect 329196 452956 329248 453008
rect 329840 452956 329892 453008
rect 330668 452956 330720 453008
rect 330760 452956 330812 453008
rect 418804 452956 418856 453008
rect 188068 452888 188120 452940
rect 261760 452888 261812 452940
rect 291936 452888 291988 452940
rect 391204 452888 391256 452940
rect 188528 452820 188580 452872
rect 265808 452820 265860 452872
rect 298192 452820 298244 452872
rect 402428 452820 402480 452872
rect 185492 452752 185544 452804
rect 262220 452752 262272 452804
rect 283472 452752 283524 452804
rect 392584 452752 392636 452804
rect 185584 452684 185636 452736
rect 263968 452684 264020 452736
rect 279056 452684 279108 452736
rect 390100 452684 390152 452736
rect 191564 452616 191616 452668
rect 270960 452616 271012 452668
rect 325792 452616 325844 452668
rect 330760 452616 330812 452668
rect 371240 452616 371292 452668
rect 372252 452616 372304 452668
rect 376760 452616 376812 452668
rect 377404 452616 377456 452668
rect 378140 452616 378192 452668
rect 378876 452616 378928 452668
rect 386144 452616 386196 452668
rect 390652 452616 390704 452668
rect 235264 452548 235316 452600
rect 236368 452548 236420 452600
rect 280804 452548 280856 452600
rect 282000 452548 282052 452600
rect 307024 452548 307076 452600
rect 308036 452548 308088 452600
rect 308128 452548 308180 452600
rect 309048 452548 309100 452600
rect 369860 452548 369912 452600
rect 378692 452548 378744 452600
rect 228364 452480 228416 452532
rect 237104 452480 237156 452532
rect 287152 452480 287204 452532
rect 288348 452480 288400 452532
rect 387616 452480 387668 452532
rect 228456 452412 228508 452464
rect 237840 452412 237892 452464
rect 228732 452344 228784 452396
rect 259184 452344 259236 452396
rect 300032 452344 300084 452396
rect 300768 452344 300820 452396
rect 390192 452412 390244 452464
rect 377312 452344 377364 452396
rect 418896 452344 418948 452396
rect 203616 452276 203668 452328
rect 214564 452276 214616 452328
rect 232596 452276 232648 452328
rect 252928 452276 252980 452328
rect 308496 452276 308548 452328
rect 417424 452276 417476 452328
rect 203984 452208 204036 452260
rect 214472 452208 214524 452260
rect 228548 452208 228600 452260
rect 258080 452208 258132 452260
rect 364432 452208 364484 452260
rect 3516 452140 3568 452192
rect 234988 452140 235040 452192
rect 235356 452140 235408 452192
rect 277216 452140 277268 452192
rect 317696 452140 317748 452192
rect 370320 452208 370372 452260
rect 378968 452208 379020 452260
rect 191380 452072 191432 452124
rect 226800 452072 226852 452124
rect 232688 452072 232740 452124
rect 275008 452072 275060 452124
rect 310704 452072 310756 452124
rect 377864 452140 377916 452192
rect 190920 452004 190972 452056
rect 228364 452004 228416 452056
rect 228640 452004 228692 452056
rect 189632 451936 189684 451988
rect 228916 451936 228968 451988
rect 232872 452004 232924 452056
rect 276480 452004 276532 452056
rect 306656 452004 306708 452056
rect 369860 452004 369912 452056
rect 378784 452072 378836 452124
rect 379060 452004 379112 452056
rect 255504 451936 255556 451988
rect 257344 451936 257396 451988
rect 366272 451936 366324 451988
rect 367376 451936 367428 451988
rect 191288 451868 191340 451920
rect 231952 451868 232004 451920
rect 232504 451868 232556 451920
rect 254400 451868 254452 451920
rect 255872 451868 255924 451920
rect 369124 451868 369176 451920
rect 379152 451868 379204 451920
rect 380256 451868 380308 451920
rect 388628 451868 388680 451920
rect 177304 451800 177356 451852
rect 227168 451800 227220 451852
rect 378140 451800 378192 451852
rect 389916 451800 389968 451852
rect 185676 451732 185728 451784
rect 275744 451732 275796 451784
rect 322480 451732 322532 451784
rect 388812 451732 388864 451784
rect 48964 451664 49016 451716
rect 232688 451664 232740 451716
rect 296720 451664 296772 451716
rect 372528 451664 372580 451716
rect 372896 451664 372948 451716
rect 416044 451664 416096 451716
rect 214564 451596 214616 451648
rect 387708 451596 387760 451648
rect 188896 451528 188948 451580
rect 195520 451528 195572 451580
rect 214472 451528 214524 451580
rect 388904 451528 388956 451580
rect 19708 451460 19760 451512
rect 232320 451460 232372 451512
rect 383200 451460 383252 451512
rect 413284 451460 413336 451512
rect 19984 451392 20036 451444
rect 234528 451392 234580 451444
rect 3608 451324 3660 451376
rect 231216 451324 231268 451376
rect 308128 451324 308180 451376
rect 383660 451324 383712 451376
rect 188620 451256 188672 451308
rect 188896 451256 188948 451308
rect 205916 451256 205968 451308
rect 206100 451256 206152 451308
rect 204260 451188 204312 451240
rect 226432 451256 226484 451308
rect 381728 451256 381780 451308
rect 389824 451392 389876 451444
rect 384672 451324 384724 451376
rect 390008 451324 390060 451376
rect 385408 451256 385460 451308
rect 388076 451256 388128 451308
rect 242900 451052 242952 451104
rect 243360 451052 243412 451104
rect 219624 450984 219676 451036
rect 219808 450984 219860 451036
rect 158076 450916 158128 450968
rect 345664 450916 345716 450968
rect 156604 450848 156656 450900
rect 339776 450848 339828 450900
rect 341984 450848 342036 450900
rect 416320 450848 416372 450900
rect 156696 450780 156748 450832
rect 351552 450780 351604 450832
rect 191104 450712 191156 450764
rect 226064 450712 226116 450764
rect 374368 450712 374420 450764
rect 411076 450712 411128 450764
rect 188252 450644 188304 450696
rect 227904 450644 227956 450696
rect 371424 450644 371476 450696
rect 410984 450644 411036 450696
rect 182824 450576 182876 450628
rect 230848 450576 230900 450628
rect 368480 450576 368532 450628
rect 410892 450576 410944 450628
rect 3700 450508 3752 450560
rect 204260 450508 204312 450560
rect 219440 450508 219492 450560
rect 219900 450508 219952 450560
rect 220912 450508 220964 450560
rect 221372 450508 221424 450560
rect 356704 450508 356756 450560
rect 189816 450440 189868 450492
rect 269856 450440 269908 450492
rect 358912 450440 358964 450492
rect 359096 450440 359148 450492
rect 359648 450508 359700 450560
rect 410800 450508 410852 450560
rect 413468 450440 413520 450492
rect 187424 450372 187476 450424
rect 269488 450372 269540 450424
rect 276112 450372 276164 450424
rect 276572 450372 276624 450424
rect 285772 450372 285824 450424
rect 286048 450372 286100 450424
rect 353760 450372 353812 450424
rect 413560 450372 413612 450424
rect 184112 450304 184164 450356
rect 288624 450304 288676 450356
rect 302240 450304 302292 450356
rect 302608 450304 302660 450356
rect 350816 450304 350868 450356
rect 413652 450304 413704 450356
rect 191196 450236 191248 450288
rect 305552 450236 305604 450288
rect 347872 450236 347924 450288
rect 413744 450236 413796 450288
rect 182088 450168 182140 450220
rect 297456 450168 297508 450220
rect 329104 450168 329156 450220
rect 418988 450168 419040 450220
rect 212540 450100 212592 450152
rect 212908 450100 212960 450152
rect 215300 450100 215352 450152
rect 216220 450100 216272 450152
rect 216680 450100 216732 450152
rect 217324 450100 217376 450152
rect 218152 450100 218204 450152
rect 218796 450100 218848 450152
rect 219532 450100 219584 450152
rect 220268 450100 220320 450152
rect 221004 450100 221056 450152
rect 221740 450100 221792 450152
rect 222200 450100 222252 450152
rect 223212 450100 223264 450152
rect 259460 450100 259512 450152
rect 260012 450100 260064 450152
rect 332416 450100 332468 450152
rect 416136 450100 416188 450152
rect 212632 450032 212684 450084
rect 213276 450032 213328 450084
rect 216772 450032 216824 450084
rect 217692 450032 217744 450084
rect 220820 450032 220872 450084
rect 221188 450032 221240 450084
rect 335636 450032 335688 450084
rect 416412 450032 416464 450084
rect 158168 449964 158220 450016
rect 336280 449964 336332 450016
rect 338948 449964 339000 450016
rect 416228 449964 416280 450016
rect 191840 449896 191892 449948
rect 225512 449896 225564 449948
rect 314660 449896 314712 449948
rect 314936 449896 314988 449948
rect 365720 449896 365772 449948
rect 388536 449896 388588 449948
rect 3332 449828 3384 449880
rect 193864 449828 193916 449880
rect 387708 449760 387760 449812
rect 388996 449760 389048 449812
rect 349620 449692 349672 449744
rect 405556 449692 405608 449744
rect 190184 449624 190236 449676
rect 263508 449624 263560 449676
rect 312820 449624 312872 449676
rect 407672 449624 407724 449676
rect 189908 449556 189960 449608
rect 267464 449556 267516 449608
rect 189724 449488 189776 449540
rect 268568 449556 268620 449608
rect 309048 449556 309100 449608
rect 408224 449556 408276 449608
rect 388996 449488 389048 449540
rect 580908 449488 580960 449540
rect 188436 447924 188488 447976
rect 188620 447924 188672 447976
rect 188068 446428 188120 446480
rect 188436 446428 188488 446480
rect 388904 442212 388956 442264
rect 580816 442212 580868 442264
rect 390376 422900 390428 422952
rect 580816 422900 580868 422952
rect 394148 419432 394200 419484
rect 580172 419432 580224 419484
rect 3332 398760 3384 398812
rect 190828 398760 190880 398812
rect 189540 397400 189592 397452
rect 190828 397400 190880 397452
rect 390284 379448 390336 379500
rect 580172 379448 580224 379500
rect 3056 372512 3108 372564
rect 190828 372512 190880 372564
rect 399760 365644 399812 365696
rect 580172 365644 580224 365696
rect 3332 358708 3384 358760
rect 184020 358708 184072 358760
rect 395436 353200 395488 353252
rect 580172 353200 580224 353252
rect 3332 346332 3384 346384
rect 177304 346332 177356 346384
rect 391296 325592 391348 325644
rect 580172 325592 580224 325644
rect 2964 320084 3016 320136
rect 188252 320084 188304 320136
rect 403624 313216 403676 313268
rect 580172 313216 580224 313268
rect 3332 306280 3384 306332
rect 190920 306280 190972 306332
rect 2872 293904 2924 293956
rect 181352 293904 181404 293956
rect 395344 273164 395396 273216
rect 580172 273164 580224 273216
rect 3240 267656 3292 267708
rect 189632 267656 189684 267708
rect 396724 259360 396776 259412
rect 579804 259360 579856 259412
rect 3332 255212 3384 255264
rect 190920 255212 190972 255264
rect 186872 250452 186924 250504
rect 218704 250452 218756 250504
rect 378232 249704 378284 249756
rect 386420 249704 386472 249756
rect 386420 248412 386472 248464
rect 389364 248412 389416 248464
rect 216404 248344 216456 248396
rect 236092 248344 236144 248396
rect 313372 248344 313424 248396
rect 358360 248344 358412 248396
rect 383752 248344 383804 248396
rect 389180 248344 389232 248396
rect 217600 248276 217652 248328
rect 237472 248276 237524 248328
rect 314752 248276 314804 248328
rect 360936 248276 360988 248328
rect 385132 248276 385184 248328
rect 389272 248276 389324 248328
rect 217508 248208 217560 248260
rect 238852 248208 238904 248260
rect 316132 248208 316184 248260
rect 363604 248208 363656 248260
rect 382372 248208 382424 248260
rect 388168 248208 388220 248260
rect 217968 248140 218020 248192
rect 240232 248140 240284 248192
rect 311992 248140 312044 248192
rect 359556 248140 359608 248192
rect 379612 248140 379664 248192
rect 391940 248140 391992 248192
rect 182916 248072 182968 248124
rect 201592 248072 201644 248124
rect 217876 248072 217928 248124
rect 241612 248072 241664 248124
rect 276112 248072 276164 248124
rect 357532 248072 357584 248124
rect 380992 248072 381044 248124
rect 390560 248072 390612 248124
rect 181352 248004 181404 248056
rect 200212 248004 200264 248056
rect 217784 248004 217836 248056
rect 242992 248004 243044 248056
rect 305092 248004 305144 248056
rect 402980 248004 403032 248056
rect 179236 247936 179288 247988
rect 204352 247936 204404 247988
rect 219348 247936 219400 247988
rect 245752 247936 245804 247988
rect 299572 247936 299624 247988
rect 304264 247936 304316 247988
rect 306472 247936 306524 247988
rect 407120 247936 407172 247988
rect 174544 247868 174596 247920
rect 207112 247868 207164 247920
rect 217692 247868 217744 247920
rect 244372 247868 244424 247920
rect 307852 247868 307904 247920
rect 409880 247868 409932 247920
rect 175832 247800 175884 247852
rect 208492 247800 208544 247852
rect 216588 247800 216640 247852
rect 248512 247800 248564 247852
rect 309232 247800 309284 247852
rect 414020 247800 414072 247852
rect 1400 247732 1452 247784
rect 193312 247732 193364 247784
rect 215208 247732 215260 247784
rect 247132 247732 247184 247784
rect 267832 247732 267884 247784
rect 356612 247732 356664 247784
rect 387892 247732 387944 247784
rect 558920 247732 558972 247784
rect 20 247664 72 247716
rect 191932 247664 191984 247716
rect 216496 247664 216548 247716
rect 249892 247664 249944 247716
rect 271972 247664 272024 247716
rect 361672 247664 361724 247716
rect 376852 247664 376904 247716
rect 582380 247664 582432 247716
rect 211252 247596 211304 247648
rect 230572 247596 230624 247648
rect 320272 247596 320324 247648
rect 358176 247596 358228 247648
rect 217416 247528 217468 247580
rect 234712 247528 234764 247580
rect 331312 247528 331364 247580
rect 359464 247528 359516 247580
rect 215300 247460 215352 247512
rect 231952 247460 232004 247512
rect 338212 247460 338264 247512
rect 356704 247460 356756 247512
rect 291292 247120 291344 247172
rect 293224 247120 293276 247172
rect 298192 247120 298244 247172
rect 302884 247120 302936 247172
rect 195244 247052 195296 247104
rect 196072 247052 196124 247104
rect 231124 247052 231176 247104
rect 233332 247052 233384 247104
rect 289912 247052 289964 247104
rect 291844 247052 291896 247104
rect 294052 247052 294104 247104
rect 295984 247052 296036 247104
rect 296812 247052 296864 247104
rect 298744 247052 298796 247104
rect 300952 247052 301004 247104
rect 305644 247052 305696 247104
rect 165620 246304 165672 246356
rect 212632 246304 212684 246356
rect 292672 246304 292724 246356
rect 371240 246304 371292 246356
rect 386420 246304 386472 246356
rect 415400 246304 415452 246356
rect 387064 245624 387116 245676
rect 387892 245624 387944 245676
rect 392676 245556 392728 245608
rect 580172 245556 580224 245608
rect 161480 244876 161532 244928
rect 211160 244876 211212 244928
rect 325792 244876 325844 244928
rect 411904 244876 411956 244928
rect 332692 243584 332744 243636
rect 381544 243584 381596 243636
rect 172520 243516 172572 243568
rect 215392 243516 215444 243568
rect 368572 243516 368624 243568
rect 565820 243516 565872 243568
rect 176660 242156 176712 242208
rect 216772 242156 216824 242208
rect 371332 242156 371384 242208
rect 565084 242156 565136 242208
rect 3240 241408 3292 241460
rect 185400 241408 185452 241460
rect 295340 239436 295392 239488
rect 378140 239436 378192 239488
rect 179420 239368 179472 239420
rect 218060 239368 218112 239420
rect 372620 239368 372672 239420
rect 569224 239368 569276 239420
rect 293224 236648 293276 236700
rect 367192 236648 367244 236700
rect 374000 236648 374052 236700
rect 578884 236648 578936 236700
rect 328460 233860 328512 233912
rect 408408 233860 408460 233912
rect 298744 232500 298796 232552
rect 382280 232500 382332 232552
rect 302884 229712 302936 229764
rect 385040 229712 385092 229764
rect 3792 217268 3844 217320
rect 191288 217268 191340 217320
rect 3332 215228 3384 215280
rect 187332 215228 187384 215280
rect 394056 206932 394108 206984
rect 579804 206932 579856 206984
rect 3332 202784 3384 202836
rect 182824 202784 182876 202836
rect 375380 199384 375432 199436
rect 562416 199384 562468 199436
rect 369860 197956 369912 198008
rect 569960 197956 570012 198008
rect 150992 195984 151044 196036
rect 157340 195984 157392 196036
rect 551008 195984 551060 196036
rect 557540 195984 557592 196036
rect 18420 195508 18472 195560
rect 34520 195508 34572 195560
rect 17132 195440 17184 195492
rect 52460 195440 52512 195492
rect 18696 195372 18748 195424
rect 66260 195372 66312 195424
rect 19616 195304 19668 195356
rect 80152 195304 80204 195356
rect 18512 195236 18564 195288
rect 80060 195236 80112 195288
rect 3700 193808 3752 193860
rect 48964 193808 49016 193860
rect 562324 193128 562376 193180
rect 579620 193128 579672 193180
rect 3332 188980 3384 189032
rect 18604 188980 18656 189032
rect 310520 180072 310572 180124
rect 416504 180072 416556 180124
rect 570604 166948 570656 167000
rect 580172 166948 580224 167000
rect 573364 153144 573416 153196
rect 580172 153144 580224 153196
rect 405648 146888 405700 146940
rect 416780 146888 416832 146940
rect 413928 144848 413980 144900
rect 417148 144848 417200 144900
rect 411168 141380 411220 141432
rect 416780 141380 416832 141432
rect 409788 140020 409840 140072
rect 416780 140020 416832 140072
rect 15936 138252 15988 138304
rect 17868 138252 17920 138304
rect 3056 137912 3108 137964
rect 10324 137912 10376 137964
rect 417148 137300 417200 137352
rect 417608 137300 417660 137352
rect 333980 129004 334032 129056
rect 406384 129004 406436 129056
rect 327080 127576 327132 127628
rect 413836 127576 413888 127628
rect 566464 126896 566516 126948
rect 580172 126896 580224 126948
rect 324320 126216 324372 126268
rect 416596 126216 416648 126268
rect 322940 124856 322992 124908
rect 414664 124856 414716 124908
rect 321560 123428 321612 123480
rect 415952 123428 416004 123480
rect 291844 122068 291896 122120
rect 364432 122068 364484 122120
rect 287060 120708 287112 120760
rect 357624 120708 357676 120760
rect 417792 120164 417844 120216
rect 419264 120164 419316 120216
rect 351184 117920 351236 117972
rect 415400 117920 415452 117972
rect 417792 117920 417844 117972
rect 305644 115200 305696 115252
rect 391940 115200 391992 115252
rect 304264 113772 304316 113824
rect 389180 113772 389232 113824
rect 571984 113092 572036 113144
rect 579988 113092 580040 113144
rect 295984 112548 296036 112600
rect 374000 112548 374052 112600
rect 303620 112480 303672 112532
rect 398840 112480 398892 112532
rect 318800 112412 318852 112464
rect 419080 112412 419132 112464
rect 3332 111732 3384 111784
rect 19708 111732 19760 111784
rect 288440 111188 288492 111240
rect 360292 111188 360344 111240
rect 302240 111120 302292 111172
rect 396080 111120 396132 111172
rect 317420 111052 317472 111104
rect 418528 111052 418580 111104
rect 417976 109692 418028 109744
rect 451280 109692 451332 109744
rect 452476 109692 452528 109744
rect 418988 109624 419040 109676
rect 480904 109624 480956 109676
rect 416136 109556 416188 109608
rect 483480 109556 483532 109608
rect 416412 109488 416464 109540
rect 485964 109488 486016 109540
rect 416228 109420 416280 109472
rect 488264 109420 488316 109472
rect 416320 109352 416372 109404
rect 491024 109352 491076 109404
rect 413376 109284 413428 109336
rect 493416 109284 493468 109336
rect 413744 109216 413796 109268
rect 495900 109216 495952 109268
rect 413652 109148 413704 109200
rect 498476 109148 498528 109200
rect 388812 109080 388864 109132
rect 476120 109080 476172 109132
rect 410708 109012 410760 109064
rect 508504 109012 508556 109064
rect 113456 108944 113508 108996
rect 184388 108944 184440 108996
rect 111064 108876 111116 108928
rect 184296 108876 184348 108928
rect 108580 108808 108632 108860
rect 184480 108808 184532 108860
rect 413560 108808 413612 108860
rect 500960 108808 501012 108860
rect 106004 108740 106056 108792
rect 184204 108740 184256 108792
rect 413468 108740 413520 108792
rect 503444 108740 503496 108792
rect 100944 108672 100996 108724
rect 184664 108672 184716 108724
rect 410800 108672 410852 108724
rect 505928 108672 505980 108724
rect 68376 108604 68428 108656
rect 181904 108604 181956 108656
rect 412548 108604 412600 108656
rect 416136 108604 416188 108656
rect 418896 108604 418948 108656
rect 520924 108604 520976 108656
rect 61108 108536 61160 108588
rect 181720 108536 181772 108588
rect 410892 108536 410944 108588
rect 513380 108536 513432 108588
rect 56048 108468 56100 108520
rect 181996 108468 182048 108520
rect 410984 108468 411036 108520
rect 515864 108468 515916 108520
rect 53656 108400 53708 108452
rect 184112 108400 184164 108452
rect 411076 108400 411128 108452
rect 518440 108400 518492 108452
rect 50804 108332 50856 108384
rect 184572 108332 184624 108384
rect 413284 108332 413336 108384
rect 525892 108332 525944 108384
rect 48320 108264 48372 108316
rect 187240 108264 187292 108316
rect 285680 108264 285732 108316
rect 358820 108264 358872 108316
rect 388628 108264 388680 108316
rect 523316 108264 523368 108316
rect 414388 108196 414440 108248
rect 414848 108196 414900 108248
rect 415124 108128 415176 108180
rect 416412 108128 416464 108180
rect 18420 108060 18472 108112
rect 19248 108060 19300 108112
rect 19524 107992 19576 108044
rect 19800 107992 19852 108044
rect 414572 107992 414624 108044
rect 415216 107992 415268 108044
rect 457996 107992 458048 108044
rect 418068 107924 418120 107976
rect 418436 107924 418488 107976
rect 452568 107924 452620 107976
rect 418344 107856 418396 107908
rect 419264 107856 419316 107908
rect 456984 107856 457036 107908
rect 19248 107788 19300 107840
rect 16488 107720 16540 107772
rect 19616 107720 19668 107772
rect 18696 107584 18748 107636
rect 19432 107584 19484 107636
rect 416412 107788 416464 107840
rect 455788 107788 455840 107840
rect 416136 107720 416188 107772
rect 458180 107720 458232 107772
rect 50160 107652 50212 107704
rect 416320 107652 416372 107704
rect 418160 107652 418212 107704
rect 418896 107652 418948 107704
rect 456984 107652 457036 107704
rect 59636 107584 59688 107636
rect 63592 107584 63644 107636
rect 191196 107584 191248 107636
rect 392584 107584 392636 107636
rect 450636 107584 450688 107636
rect 458180 107584 458232 107636
rect 459468 107584 459520 107636
rect 19064 107516 19116 107568
rect 36912 107516 36964 107568
rect 50160 107516 50212 107568
rect 68652 107516 68704 107568
rect 73712 107516 73764 107568
rect 186964 107516 187016 107568
rect 408132 107516 408184 107568
rect 458364 107516 458416 107568
rect 475660 107584 475712 107636
rect 478052 107516 478104 107568
rect 18512 107448 18564 107500
rect 19616 107448 19668 107500
rect 16120 107380 16172 107432
rect 18788 107380 18840 107432
rect 18972 107380 19024 107432
rect 35900 107380 35952 107432
rect 19156 107312 19208 107364
rect 38108 107312 38160 107364
rect 18880 107244 18932 107296
rect 39580 107244 39632 107296
rect 19708 107176 19760 107228
rect 43168 107448 43220 107500
rect 61660 107448 61712 107500
rect 61752 107448 61804 107500
rect 75644 107448 75696 107500
rect 76104 107448 76156 107500
rect 187148 107448 187200 107500
rect 408040 107448 408092 107500
rect 455972 107448 456024 107500
rect 52276 107380 52328 107432
rect 69756 107380 69808 107432
rect 78496 107380 78548 107432
rect 187056 107380 187108 107432
rect 417884 107380 417936 107432
rect 419264 107380 419316 107432
rect 455788 107380 455840 107432
rect 474372 107448 474424 107500
rect 44364 107312 44416 107364
rect 45376 107312 45428 107364
rect 63868 107312 63920 107364
rect 86040 107312 86092 107364
rect 158168 107312 158220 107364
rect 418896 107312 418948 107364
rect 46572 107244 46624 107296
rect 65156 107244 65208 107296
rect 88248 107244 88300 107296
rect 156604 107244 156656 107296
rect 19524 107108 19576 107160
rect 44272 107176 44324 107228
rect 48780 107176 48832 107228
rect 67640 107176 67692 107228
rect 93584 107176 93636 107228
rect 158076 107176 158128 107228
rect 418712 107176 418764 107228
rect 436100 107176 436152 107228
rect 452568 107312 452620 107364
rect 471152 107380 471204 107432
rect 452476 107244 452528 107296
rect 469772 107244 469824 107296
rect 459560 107176 459612 107228
rect 44180 107108 44232 107160
rect 47584 107108 47636 107160
rect 66260 107108 66312 107160
rect 121000 107108 121052 107160
rect 181812 107108 181864 107160
rect 419816 107108 419868 107160
rect 438124 107108 438176 107160
rect 444288 107108 444340 107160
rect 461676 107108 461728 107160
rect 17132 107040 17184 107092
rect 52368 107040 52420 107092
rect 15568 106972 15620 107024
rect 16212 106972 16264 107024
rect 51264 106972 51316 107024
rect 52276 106972 52328 107024
rect 59360 107040 59412 107092
rect 60556 107040 60608 107092
rect 79140 107040 79192 107092
rect 123392 107040 123444 107092
rect 181628 107040 181680 107092
rect 419724 107040 419776 107092
rect 439596 107040 439648 107092
rect 71228 106972 71280 107024
rect 98552 106972 98604 107024
rect 156696 106972 156748 107024
rect 339500 106972 339552 107024
rect 359648 106972 359700 107024
rect 415124 106972 415176 107024
rect 444196 107040 444248 107092
rect 462780 107040 462832 107092
rect 15016 106904 15068 106956
rect 53472 106904 53524 106956
rect 72148 106904 72200 106956
rect 335360 106904 335412 106956
rect 418896 106904 418948 106956
rect 419908 106904 419960 106956
rect 454592 106972 454644 107024
rect 473360 106972 473412 107024
rect 459560 106904 459612 106956
rect 460664 106904 460716 106956
rect 479156 106904 479208 106956
rect 59636 106836 59688 106888
rect 77668 106836 77720 106888
rect 418988 106836 419040 106888
rect 419356 106836 419408 106888
rect 437020 106836 437072 106888
rect 44272 106768 44324 106820
rect 62580 106768 62632 106820
rect 410616 106768 410668 106820
rect 453580 106768 453632 106820
rect 448520 106632 448572 106684
rect 467012 106632 467064 106684
rect 447140 106564 447192 106616
rect 465724 106564 465776 106616
rect 19800 106496 19852 106548
rect 40500 106496 40552 106548
rect 42800 106496 42852 106548
rect 48780 106496 48832 106548
rect 449900 106496 449952 106548
rect 468668 106496 468720 106548
rect 18328 106428 18380 106480
rect 18788 106428 18840 106480
rect 44364 106428 44416 106480
rect 55772 106428 55824 106480
rect 74356 106428 74408 106480
rect 418068 106428 418120 106480
rect 440516 106428 440568 106480
rect 445668 106428 445720 106480
rect 463884 106428 463936 106480
rect 19432 106360 19484 106412
rect 46572 106360 46624 106412
rect 55312 106360 55364 106412
rect 73252 106360 73304 106412
rect 417056 106360 417108 106412
rect 441620 106360 441672 106412
rect 446404 106360 446456 106412
rect 465172 106360 465224 106412
rect 19616 106292 19668 106344
rect 59360 106292 59412 106344
rect 419264 106292 419316 106344
rect 443092 106292 443144 106344
rect 444288 106292 444340 106344
rect 453948 106292 454000 106344
rect 472072 106292 472124 106344
rect 17224 106224 17276 106276
rect 150808 106224 150860 106276
rect 157340 106224 157392 106276
rect 351184 106224 351236 106276
rect 415032 106224 415084 106276
rect 416228 106224 416280 106276
rect 417792 106224 417844 106276
rect 550732 106224 550784 106276
rect 557540 106224 557592 106276
rect 14832 106156 14884 106208
rect 15108 106156 15160 106208
rect 44180 106156 44232 106208
rect 414480 106156 414532 106208
rect 415308 106156 415360 106208
rect 417700 106156 417752 106208
rect 418620 106156 418672 106208
rect 420000 106156 420052 106208
rect 453948 106156 454000 106208
rect 16028 106088 16080 106140
rect 16396 106088 16448 106140
rect 42800 106088 42852 106140
rect 447140 106088 447192 106140
rect 414756 106020 414808 106072
rect 446404 106020 446456 106072
rect 219164 105952 219216 106004
rect 251180 105952 251232 106004
rect 280160 105952 280212 106004
rect 357256 105952 357308 106004
rect 414572 105952 414624 106004
rect 445668 105952 445720 106004
rect 219992 105884 220044 105936
rect 252560 105884 252612 105936
rect 278780 105884 278832 105936
rect 357900 105884 357952 105936
rect 219256 105816 219308 105868
rect 255320 105816 255372 105868
rect 277400 105816 277452 105868
rect 357716 105816 357768 105868
rect 217232 105748 217284 105800
rect 259460 105748 259512 105800
rect 274640 105748 274692 105800
rect 357808 105748 357860 105800
rect 15660 105680 15712 105732
rect 18604 105680 18656 105732
rect 55312 105680 55364 105732
rect 216220 105680 216272 105732
rect 262220 105680 262272 105732
rect 273260 105680 273312 105732
rect 357072 105680 357124 105732
rect 15844 105612 15896 105664
rect 18512 105612 18564 105664
rect 55772 105612 55824 105664
rect 216312 105612 216364 105664
rect 263600 105612 263652 105664
rect 270500 105612 270552 105664
rect 358912 105612 358964 105664
rect 418620 105612 418672 105664
rect 449900 105612 449952 105664
rect 16304 105544 16356 105596
rect 18696 105544 18748 105596
rect 57060 105544 57112 105596
rect 218980 105544 219032 105596
rect 266360 105544 266412 105596
rect 269120 105544 269172 105596
rect 359004 105544 359056 105596
rect 414388 105544 414440 105596
rect 414756 105544 414808 105596
rect 416228 105544 416280 105596
rect 448520 105544 448572 105596
rect 17040 104796 17092 104848
rect 390652 104796 390704 104848
rect 417148 104796 417200 104848
rect 417424 104796 417476 104848
rect 219900 104728 219952 104780
rect 222844 104728 222896 104780
rect 219716 104660 219768 104712
rect 228364 104660 228416 104712
rect 351920 104592 351972 104644
rect 411996 104592 412048 104644
rect 350540 104524 350592 104576
rect 414940 104524 414992 104576
rect 219808 104456 219860 104508
rect 223028 104456 223080 104508
rect 349160 104456 349212 104508
rect 414756 104456 414808 104508
rect 346400 104388 346452 104440
rect 414848 104388 414900 104440
rect 219072 104320 219124 104372
rect 225604 104320 225656 104372
rect 284300 104320 284352 104372
rect 359096 104320 359148 104372
rect 282920 104252 282972 104304
rect 359280 104252 359332 104304
rect 217140 104184 217192 104236
rect 225788 104184 225840 104236
rect 281540 104184 281592 104236
rect 359188 104184 359240 104236
rect 218060 104116 218112 104168
rect 231124 104116 231176 104168
rect 329840 104116 329892 104168
rect 418804 104116 418856 104168
rect 216128 103504 216180 103556
rect 359740 103504 359792 103556
rect 183560 102756 183612 102808
rect 219440 102756 219492 102808
rect 360108 99288 360160 99340
rect 387064 99288 387116 99340
rect 356980 98744 357032 98796
rect 158904 98608 158956 98660
rect 170496 98608 170548 98660
rect 357164 98608 357216 98660
rect 356980 98540 357032 98592
rect 357164 98404 357216 98456
rect 3332 71680 3384 71732
rect 14556 71680 14608 71732
rect 3332 59304 3384 59356
rect 14464 59304 14516 59356
rect 170496 57876 170548 57928
rect 216128 57876 216180 57928
rect 216680 57876 216732 57928
rect 191564 56516 191616 56568
rect 216680 56516 216732 56568
rect 189816 53728 189868 53780
rect 216680 53728 216732 53780
rect 189724 53660 189776 53712
rect 216772 53660 216824 53712
rect 189908 52368 189960 52420
rect 216772 52368 216824 52420
rect 190000 51008 190052 51060
rect 216680 51008 216732 51060
rect 190092 48220 190144 48272
rect 216680 48220 216732 48272
rect 558184 46860 558236 46912
rect 580172 46860 580224 46912
rect 3332 45500 3384 45552
rect 7564 45500 7616 45552
rect 3332 33056 3384 33108
rect 19984 33056 20036 33108
rect 391204 28908 391256 28960
rect 416780 28908 416832 28960
rect 371148 28228 371200 28280
rect 416872 28228 416924 28280
rect 418712 22584 418764 22636
rect 419172 22584 419224 22636
rect 418436 22380 418488 22432
rect 418620 22380 418672 22432
rect 217324 20000 217376 20052
rect 371148 20000 371200 20052
rect 416320 19728 416372 19780
rect 460664 19728 460716 19780
rect 405464 19660 405516 19712
rect 488264 19660 488316 19712
rect 405096 19592 405148 19644
rect 491024 19592 491076 19644
rect 405280 19524 405332 19576
rect 493416 19524 493468 19576
rect 405556 19456 405608 19508
rect 495900 19456 495952 19508
rect 17132 19388 17184 19440
rect 52368 19388 52420 19440
rect 402704 19388 402756 19440
rect 500960 19388 501012 19440
rect 15016 19320 15068 19372
rect 53472 19320 53524 19372
rect 188988 19320 189040 19372
rect 285956 19320 286008 19372
rect 402796 19320 402848 19372
rect 503536 19320 503588 19372
rect 103704 19252 103756 19304
rect 176200 19252 176252 19304
rect 188804 19252 188856 19304
rect 244280 19252 244332 19304
rect 415308 19252 415360 19304
rect 447600 19252 447652 19304
rect 100944 19184 100996 19236
rect 176292 19184 176344 19236
rect 190276 19184 190328 19236
rect 246396 19184 246448 19236
rect 416228 19184 416280 19236
rect 448704 19184 448756 19236
rect 95976 19116 96028 19168
rect 176568 19116 176620 19168
rect 188528 19116 188580 19168
rect 245292 19116 245344 19168
rect 416412 19116 416464 19168
rect 455972 19116 456024 19168
rect 91008 19048 91060 19100
rect 178592 19048 178644 19100
rect 188620 19048 188672 19100
rect 248236 19048 248288 19100
rect 399484 19048 399536 19100
rect 468300 19048 468352 19100
rect 86040 18980 86092 19032
rect 179144 18980 179196 19032
rect 191748 18980 191800 19032
rect 250076 18980 250128 19032
rect 399576 18980 399628 19032
rect 470876 18980 470928 19032
rect 81072 18912 81124 18964
rect 179328 18912 179380 18964
rect 187516 18912 187568 18964
rect 247500 18912 247552 18964
rect 416044 18912 416096 18964
rect 515772 18912 515824 18964
rect 76104 18844 76156 18896
rect 179052 18844 179104 18896
rect 190184 18844 190236 18896
rect 250628 18844 250680 18896
rect 402612 18844 402664 18896
rect 505836 18844 505888 18896
rect 18420 18776 18472 18828
rect 58164 18776 58216 18828
rect 73712 18776 73764 18828
rect 181536 18776 181588 18828
rect 190368 18776 190420 18828
rect 252284 18776 252336 18828
rect 402520 18776 402572 18828
rect 508412 18776 508464 18828
rect 56048 18708 56100 18760
rect 173624 18708 173676 18760
rect 191656 18708 191708 18760
rect 253572 18708 253624 18760
rect 389916 18708 389968 18760
rect 498476 18708 498528 18760
rect 53656 18640 53708 18692
rect 173808 18640 173860 18692
rect 185860 18640 185912 18692
rect 255964 18640 256016 18692
rect 389824 18640 389876 18692
rect 523316 18640 523368 18692
rect 50896 18572 50948 18624
rect 176384 18572 176436 18624
rect 185768 18572 185820 18624
rect 258356 18572 258408 18624
rect 390008 18572 390060 18624
rect 525892 18572 525944 18624
rect 106096 18504 106148 18556
rect 176476 18504 176528 18556
rect 188712 18504 188764 18556
rect 243084 18504 243136 18556
rect 418712 18504 418764 18556
rect 450084 18504 450136 18556
rect 108672 18436 108724 18488
rect 175924 18436 175976 18488
rect 188436 18436 188488 18488
rect 236000 18436 236052 18488
rect 414572 18436 414624 18488
rect 445668 18436 445720 18488
rect 113456 18368 113508 18420
rect 176108 18368 176160 18420
rect 217416 18368 217468 18420
rect 222200 18368 222252 18420
rect 415124 18368 415176 18420
rect 444288 18368 444340 18420
rect 19064 17892 19116 17944
rect 36544 17892 36596 17944
rect 62028 17892 62080 17944
rect 173348 17892 173400 17944
rect 185676 17892 185728 17944
rect 280160 17892 280212 17944
rect 402428 17892 402480 17944
rect 458364 17892 458416 17944
rect 460664 17892 460716 17944
rect 478880 17892 478932 17944
rect 19616 17824 19668 17876
rect 60464 17824 60516 17876
rect 64696 17824 64748 17876
rect 173440 17824 173492 17876
rect 187608 17824 187660 17876
rect 277400 17824 277452 17876
rect 444288 17824 444340 17876
rect 462320 17824 462372 17876
rect 18512 17756 18564 17808
rect 55956 17756 56008 17808
rect 56508 17756 56560 17808
rect 66168 17756 66220 17808
rect 173164 17756 173216 17808
rect 191472 17756 191524 17808
rect 273260 17756 273312 17808
rect 410524 17756 410576 17808
rect 455420 17756 455472 17808
rect 455972 17756 456024 17808
rect 473360 17756 473412 17808
rect 18604 17688 18656 17740
rect 53840 17688 53892 17740
rect 68928 17688 68980 17740
rect 173256 17688 173308 17740
rect 183468 17688 183520 17740
rect 264980 17688 265032 17740
rect 414480 17688 414532 17740
rect 456800 17688 456852 17740
rect 16212 17620 16264 17672
rect 51448 17620 51500 17672
rect 78588 17620 78640 17672
rect 178776 17620 178828 17672
rect 183376 17620 183428 17672
rect 263600 17620 263652 17672
rect 445668 17620 445720 17672
rect 463700 17620 463752 17672
rect 16396 17552 16448 17604
rect 48688 17552 48740 17604
rect 49608 17552 49660 17604
rect 53472 17552 53524 17604
rect 71780 17552 71832 17604
rect 191840 17552 191892 17604
rect 270500 17552 270552 17604
rect 448704 17552 448756 17604
rect 466460 17552 466512 17604
rect 15108 17484 15160 17536
rect 47584 17484 47636 17536
rect 48228 17484 48280 17536
rect 50160 17484 50212 17536
rect 67640 17484 67692 17536
rect 83832 17484 83884 17536
rect 178684 17484 178736 17536
rect 185952 17484 186004 17536
rect 260840 17484 260892 17536
rect 419264 17484 419316 17536
rect 443092 17484 443144 17536
rect 19248 17416 19300 17468
rect 60464 17416 60516 17468
rect 78680 17416 78732 17468
rect 88248 17416 88300 17468
rect 178868 17416 178920 17468
rect 184756 17416 184808 17468
rect 259552 17416 259604 17468
rect 417056 17416 417108 17468
rect 441712 17416 441764 17468
rect 19432 17348 19484 17400
rect 18328 17280 18380 17332
rect 19524 17212 19576 17264
rect 19708 17144 19760 17196
rect 18880 17076 18932 17128
rect 38660 17076 38712 17128
rect 49608 17348 49660 17400
rect 67640 17348 67692 17400
rect 69664 17348 69716 17400
rect 75920 17348 75972 17400
rect 93584 17348 93636 17400
rect 178960 17348 179012 17400
rect 186044 17348 186096 17400
rect 259460 17348 259512 17400
rect 418068 17348 418120 17400
rect 440240 17348 440292 17400
rect 450084 17484 450136 17536
rect 467840 17484 467892 17536
rect 447600 17416 447652 17468
rect 465080 17416 465132 17468
rect 459468 17348 459520 17400
rect 48228 17280 48280 17332
rect 66260 17280 66312 17332
rect 99288 17280 99340 17332
rect 176016 17280 176068 17332
rect 186136 17280 186188 17332
rect 258080 17280 258132 17332
rect 419724 17280 419776 17332
rect 438860 17280 438912 17332
rect 456800 17280 456852 17332
rect 458088 17280 458140 17332
rect 476120 17280 476172 17332
rect 46664 17212 46716 17264
rect 65064 17212 65116 17264
rect 111708 17212 111760 17264
rect 157984 17212 158036 17264
rect 184848 17212 184900 17264
rect 256700 17212 256752 17264
rect 419816 17212 419868 17264
rect 437480 17212 437532 17264
rect 45376 17144 45428 17196
rect 63500 17144 63552 17196
rect 71688 17144 71740 17196
rect 170404 17144 170456 17196
rect 186228 17144 186280 17196
rect 255320 17144 255372 17196
rect 419172 17144 419224 17196
rect 436100 17144 436152 17196
rect 44180 17076 44232 17128
rect 62120 17076 62172 17128
rect 218704 17076 218756 17128
rect 282920 17076 282972 17128
rect 418988 17076 419040 17128
rect 436284 17076 436336 17128
rect 43076 17008 43128 17060
rect 60740 17008 60792 17060
rect 191104 17008 191156 17060
rect 251180 17008 251232 17060
rect 393964 17008 394016 17060
rect 447140 17008 447192 17060
rect 51448 16940 51500 16992
rect 69020 16940 69072 16992
rect 414388 16940 414440 16992
rect 446496 16940 446548 16992
rect 465080 17212 465132 17264
rect 16488 16872 16540 16924
rect 59544 16872 59596 16924
rect 77300 16872 77352 16924
rect 418436 16872 418488 16924
rect 449900 16872 449952 16924
rect 451280 16872 451332 16924
rect 469312 16940 469364 16992
rect 469220 16872 469272 16924
rect 473452 16872 473504 16924
rect 56508 16804 56560 16856
rect 73160 16804 73212 16856
rect 457352 16804 457404 16856
rect 474740 16804 474792 16856
rect 57888 16736 57940 16788
rect 74816 16736 74868 16788
rect 451372 16736 451424 16788
rect 452292 16736 452344 16788
rect 470876 16736 470928 16788
rect 52368 16668 52420 16720
rect 70400 16668 70452 16720
rect 452660 16668 452712 16720
rect 453488 16668 453540 16720
rect 471980 16668 472032 16720
rect 125968 16532 126020 16584
rect 388076 16532 388128 16584
rect 416136 16532 416188 16584
rect 458272 16532 458324 16584
rect 477500 16600 477552 16652
rect 418344 16464 418396 16516
rect 457352 16464 457404 16516
rect 419908 16396 419960 16448
rect 454040 16396 454092 16448
rect 469220 16396 469272 16448
rect 417976 16328 418028 16380
rect 451280 16328 451332 16380
rect 420000 16260 420052 16312
rect 452660 16260 452712 16312
rect 418620 16192 418672 16244
rect 451372 16192 451424 16244
rect 359556 15920 359608 15972
rect 420920 15920 420972 15972
rect 130568 15852 130620 15904
rect 198740 15852 198792 15904
rect 363604 15852 363656 15904
rect 432052 15852 432104 15904
rect 358360 14492 358412 14544
rect 423680 14492 423732 14544
rect 126980 14424 127032 14476
rect 197452 14424 197504 14476
rect 358176 14424 358228 14476
rect 442632 14424 442684 14476
rect 362960 13064 363012 13116
rect 552664 13064 552716 13116
rect 357440 11840 357492 11892
rect 360936 11772 360988 11824
rect 428464 11772 428516 11824
rect 359464 11704 359516 11756
rect 470600 11704 470652 11756
rect 357624 11500 357676 11552
rect 128176 10276 128228 10328
rect 195244 10276 195296 10328
rect 361580 10276 361632 10328
rect 548616 10276 548668 10328
rect 360200 8916 360252 8968
rect 545488 8916 545540 8968
rect 218888 8304 218940 8356
rect 219072 8304 219124 8356
rect 357164 7624 357216 7676
rect 527824 7624 527876 7676
rect 158904 7556 158956 7608
rect 209780 7556 209832 7608
rect 218060 7556 218112 7608
rect 219256 7556 219308 7608
rect 356980 7556 357032 7608
rect 531320 7556 531372 7608
rect 216220 6332 216272 6384
rect 293684 6332 293736 6384
rect 219716 6264 219768 6316
rect 300768 6264 300820 6316
rect 216312 6196 216364 6248
rect 297272 6196 297324 6248
rect 411996 6196 412048 6248
rect 524236 6196 524288 6248
rect 169576 6128 169628 6180
rect 213920 6128 213972 6180
rect 218980 6128 219032 6180
rect 304356 6128 304408 6180
rect 357624 6128 357676 6180
rect 538404 6128 538456 6180
rect 356704 5244 356756 5296
rect 488816 5244 488868 5296
rect 360844 5176 360896 5228
rect 495900 5176 495952 5228
rect 356796 5108 356848 5160
rect 502984 5108 503036 5160
rect 358268 5040 358320 5092
rect 506480 5040 506532 5092
rect 358084 4972 358136 5024
rect 513564 4972 513616 5024
rect 364340 4904 364392 4956
rect 556160 4904 556212 4956
rect 365720 4836 365772 4888
rect 559748 4836 559800 4888
rect 125876 4768 125928 4820
rect 194600 4768 194652 4820
rect 367100 4700 367152 4752
rect 563244 4768 563296 4820
rect 217968 4088 218020 4140
rect 237012 4088 237064 4140
rect 343364 4088 343416 4140
rect 359188 4088 359240 4140
rect 414664 4088 414716 4140
rect 449808 4088 449860 4140
rect 217876 4020 217928 4072
rect 240508 4020 240560 4072
rect 339868 4020 339920 4072
rect 357072 4020 357124 4072
rect 416596 4020 416648 4072
rect 453304 4020 453356 4072
rect 217784 3952 217836 4004
rect 244096 3952 244148 4004
rect 336280 3952 336332 4004
rect 357900 3952 357952 4004
rect 411904 3952 411956 4004
rect 456892 3952 456944 4004
rect 217692 3884 217744 3936
rect 247592 3884 247644 3936
rect 332692 3884 332744 3936
rect 357716 3884 357768 3936
rect 413836 3884 413888 3936
rect 460388 3884 460440 3936
rect 155408 3816 155460 3868
rect 175832 3816 175884 3868
rect 219348 3816 219400 3868
rect 251180 3816 251232 3868
rect 329196 3816 329248 3868
rect 357440 3816 357492 3868
rect 418804 3816 418856 3868
rect 467472 3816 467524 3868
rect 151820 3748 151872 3800
rect 174544 3748 174596 3800
rect 215208 3748 215260 3800
rect 254676 3748 254728 3800
rect 325608 3748 325660 3800
rect 357808 3748 357860 3800
rect 408408 3748 408460 3800
rect 463976 3748 464028 3800
rect 144736 3680 144788 3732
rect 179236 3680 179288 3732
rect 216588 3680 216640 3732
rect 258264 3680 258316 3732
rect 322112 3680 322164 3732
rect 356888 3680 356940 3732
rect 418896 3680 418948 3732
rect 481732 3680 481784 3732
rect 137652 3612 137704 3664
rect 182916 3612 182968 3664
rect 194416 3612 194468 3664
rect 214564 3612 214616 3664
rect 216496 3612 216548 3664
rect 261760 3612 261812 3664
rect 318524 3612 318576 3664
rect 361672 3612 361724 3664
rect 406384 3612 406436 3664
rect 478144 3612 478196 3664
rect 134156 3544 134208 3596
rect 181352 3544 181404 3596
rect 190828 3544 190880 3596
rect 213184 3544 213236 3596
rect 219072 3544 219124 3596
rect 265348 3544 265400 3596
rect 315028 3544 315080 3596
rect 358912 3544 358964 3596
rect 381544 3544 381596 3596
rect 474556 3544 474608 3596
rect 565084 3544 565136 3596
rect 573916 3544 573968 3596
rect 148324 3476 148376 3528
rect 205640 3476 205692 3528
rect 219992 3476 220044 3528
rect 268844 3476 268896 3528
rect 311440 3476 311492 3528
rect 359004 3476 359056 3528
rect 398840 3476 398892 3528
rect 400128 3476 400180 3528
rect 416504 3476 416556 3528
rect 417884 3476 417936 3528
rect 141240 3408 141292 3460
rect 202880 3408 202932 3460
rect 205088 3408 205140 3460
rect 215944 3408 215996 3460
rect 219900 3408 219952 3460
rect 272432 3408 272484 3460
rect 307944 3408 307996 3460
rect 356612 3408 356664 3460
rect 359648 3408 359700 3460
rect 217508 3340 217560 3392
rect 233424 3340 233476 3392
rect 346952 3340 347004 3392
rect 359280 3340 359332 3392
rect 217600 3272 217652 3324
rect 229836 3272 229888 3324
rect 350448 3272 350500 3324
rect 359096 3272 359148 3324
rect 216404 3204 216456 3256
rect 226340 3204 226392 3256
rect 354036 3204 354088 3256
rect 358820 3204 358872 3256
rect 414848 3340 414900 3392
rect 510068 3476 510120 3528
rect 569224 3476 569276 3528
rect 577412 3476 577464 3528
rect 492312 3408 492364 3460
rect 562416 3408 562468 3460
rect 582196 3408 582248 3460
rect 415952 3136 416004 3188
rect 446220 3340 446272 3392
rect 419080 3272 419132 3324
rect 439136 3272 439188 3324
rect 418528 3204 418580 3256
rect 435548 3204 435600 3256
rect 423680 3136 423732 3188
rect 424968 3136 425020 3188
rect 578884 3068 578936 3120
rect 581000 3068 581052 3120
rect 374000 2728 374052 2780
rect 375288 2728 375340 2780
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700262 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 40512 700330 40540 703520
rect 72988 700369 73016 703520
rect 89180 700466 89208 703520
rect 105464 700534 105492 703520
rect 137848 700602 137876 703520
rect 154132 700670 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 163504 700664 163556 700670
rect 163504 700606 163556 700612
rect 137836 700596 137888 700602
rect 137836 700538 137888 700544
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 72974 700360 73030 700369
rect 40500 700324 40552 700330
rect 72974 700295 73030 700304
rect 40500 700266 40552 700272
rect 8116 700256 8168 700262
rect 8116 700198 8168 700204
rect 14464 700256 14516 700262
rect 14464 700198 14516 700204
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 10324 670744 10376 670750
rect 10324 670686 10376 670692
rect 3422 658200 3478 658209
rect 3422 658135 3424 658144
rect 3476 658135 3478 658144
rect 7564 658164 7616 658170
rect 3424 658106 3476 658112
rect 7564 658106 7616 658112
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 4804 632120 4856 632126
rect 2832 632088 2834 632097
rect 4804 632062 4856 632068
rect 2778 632023 2834 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553586 3372 553823
rect 3332 553580 3384 553586
rect 3332 553522 3384 553528
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3436 483818 3464 566879
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3424 483812 3476 483818
rect 3424 483754 3476 483760
rect 3528 480254 3556 514791
rect 3528 480226 3648 480254
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3436 462398 3464 462567
rect 3424 462392 3476 462398
rect 3424 462334 3476 462340
rect 3620 460222 3648 480226
rect 3608 460216 3660 460222
rect 3608 460158 3660 460164
rect 4816 457638 4844 632062
rect 7576 498982 7604 658106
rect 7656 553580 7708 553586
rect 7656 553522 7708 553528
rect 7564 498976 7616 498982
rect 7564 498918 7616 498924
rect 7668 458862 7696 553522
rect 10336 485178 10364 670686
rect 11704 605872 11756 605878
rect 11704 605814 11756 605820
rect 10416 579692 10468 579698
rect 10416 579634 10468 579640
rect 10324 485172 10376 485178
rect 10324 485114 10376 485120
rect 10428 461650 10456 579634
rect 11716 475522 11744 605814
rect 11796 527196 11848 527202
rect 11796 527138 11848 527144
rect 11704 475516 11756 475522
rect 11704 475458 11756 475464
rect 10416 461644 10468 461650
rect 10416 461586 10468 461592
rect 7656 458856 7708 458862
rect 7656 458798 7708 458804
rect 4804 457632 4856 457638
rect 4804 457574 4856 457580
rect 11808 456142 11836 527138
rect 14476 461718 14504 700198
rect 150990 674928 151046 674937
rect 150990 674863 150992 674872
rect 151044 674863 151046 674872
rect 157340 674892 157392 674898
rect 150992 674834 151044 674840
rect 157340 674834 157392 674840
rect 17590 626920 17646 626929
rect 17590 626855 17646 626864
rect 17222 622840 17278 622849
rect 17222 622775 17278 622784
rect 14556 618316 14608 618322
rect 14556 618258 14608 618264
rect 14464 461712 14516 461718
rect 14464 461654 14516 461660
rect 14568 457706 14596 618258
rect 16304 589280 16356 589286
rect 16304 589222 16356 589228
rect 16120 587240 16172 587246
rect 16026 587208 16082 587217
rect 16120 587182 16172 587188
rect 16026 587143 16082 587152
rect 15108 587036 15160 587042
rect 15108 586978 15160 586984
rect 15016 586900 15068 586906
rect 15016 586842 15068 586848
rect 14924 584588 14976 584594
rect 14924 584530 14976 584536
rect 14832 498228 14884 498234
rect 14832 498170 14884 498176
rect 14556 457700 14608 457706
rect 14556 457642 14608 457648
rect 11796 456136 11848 456142
rect 11796 456078 11848 456084
rect 14464 454300 14516 454306
rect 14464 454242 14516 454248
rect 10324 454232 10376 454238
rect 10324 454174 10376 454180
rect 7564 454164 7616 454170
rect 7564 454106 7616 454112
rect 3422 452296 3478 452305
rect 3422 452231 3478 452240
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3056 372564 3108 372570
rect 3056 372506 3108 372512
rect 3068 371385 3096 372506
rect 3054 371376 3110 371385
rect 3054 371311 3110 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 2964 320136 3016 320142
rect 2964 320078 3016 320084
rect 2976 319297 3004 320078
rect 2962 319288 3018 319297
rect 2962 319223 3018 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 2872 293956 2924 293962
rect 2872 293898 2924 293904
rect 2884 293185 2912 293898
rect 2870 293176 2926 293185
rect 2870 293111 2926 293120
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3332 255264 3384 255270
rect 3332 255206 3384 255212
rect 3344 254153 3372 255206
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 1400 247784 1452 247790
rect 1400 247726 1452 247732
rect 20 247716 72 247722
rect 20 247658 72 247664
rect 32 16574 60 247658
rect 32 16546 152 16574
rect 124 354 152 16546
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 247726
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3332 202836 3384 202842
rect 3332 202778 3384 202784
rect 3344 201929 3372 202778
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3332 189032 3384 189038
rect 3332 188974 3384 188980
rect 3344 188873 3372 188974
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3056 137964 3108 137970
rect 3056 137906 3108 137912
rect 3068 136785 3096 137906
rect 3054 136776 3110 136785
rect 3054 136711 3110 136720
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 3332 59356 3384 59362
rect 3332 59298 3384 59304
rect 3344 58585 3372 59298
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3332 45552 3384 45558
rect 3330 45520 3332 45529
rect 3384 45520 3386 45529
rect 3330 45455 3386 45464
rect 3332 33108 3384 33114
rect 3332 33050 3384 33056
rect 3344 32473 3372 33050
rect 3330 32464 3386 32473
rect 3330 32399 3386 32408
rect 3436 6497 3464 452231
rect 3516 452192 3568 452198
rect 3516 452134 3568 452140
rect 3528 19417 3556 452134
rect 3608 451376 3660 451382
rect 3608 451318 3660 451324
rect 3620 162897 3648 451318
rect 3700 450560 3752 450566
rect 3700 450502 3752 450508
rect 3712 410553 3740 450502
rect 3698 410544 3754 410553
rect 3698 410479 3754 410488
rect 3792 217320 3844 217326
rect 3792 217262 3844 217268
rect 3700 193860 3752 193866
rect 3700 193802 3752 193808
rect 3606 162888 3662 162897
rect 3606 162823 3662 162832
rect 3712 84697 3740 193802
rect 3804 149841 3832 217262
rect 3790 149832 3846 149841
rect 3790 149767 3846 149776
rect 3698 84688 3754 84697
rect 3698 84623 3754 84632
rect 7576 45558 7604 454106
rect 10336 137970 10364 454174
rect 10324 137964 10376 137970
rect 10324 137906 10376 137912
rect 14476 59362 14504 454242
rect 14554 449984 14610 449993
rect 14554 449919 14610 449928
rect 14568 71738 14596 449919
rect 14844 106214 14872 498170
rect 14936 497570 14964 584530
rect 15028 498506 15056 586842
rect 15016 498500 15068 498506
rect 15016 498442 15068 498448
rect 15028 498234 15056 498442
rect 15016 498228 15068 498234
rect 15016 498170 15068 498176
rect 14936 497542 15056 497570
rect 15028 497486 15056 497542
rect 15016 497480 15068 497486
rect 15016 497422 15068 497428
rect 15028 106962 15056 497422
rect 15120 496738 15148 586978
rect 15844 586696 15896 586702
rect 15844 586638 15896 586644
rect 15752 501016 15804 501022
rect 15752 500958 15804 500964
rect 15660 499656 15712 499662
rect 15660 499598 15712 499604
rect 15568 499588 15620 499594
rect 15568 499530 15620 499536
rect 15108 496732 15160 496738
rect 15108 496674 15160 496680
rect 15580 107030 15608 499530
rect 15568 107024 15620 107030
rect 15568 106966 15620 106972
rect 15016 106956 15068 106962
rect 15016 106898 15068 106904
rect 14832 106208 14884 106214
rect 14832 106150 14884 106156
rect 14556 71732 14608 71738
rect 14556 71674 14608 71680
rect 14464 59356 14516 59362
rect 14464 59298 14516 59304
rect 7564 45552 7616 45558
rect 7564 45494 7616 45500
rect 3514 19408 3570 19417
rect 15028 19378 15056 106898
rect 15108 106208 15160 106214
rect 15108 106150 15160 106156
rect 3514 19343 3570 19352
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 15120 17542 15148 106150
rect 15672 105738 15700 499598
rect 15764 458930 15792 500958
rect 15856 498302 15884 586638
rect 15934 521520 15990 521529
rect 15934 521455 15990 521464
rect 15844 498296 15896 498302
rect 15844 498238 15896 498244
rect 15752 458924 15804 458930
rect 15752 458866 15804 458872
rect 15660 105732 15712 105738
rect 15660 105674 15712 105680
rect 15856 105670 15884 498238
rect 15948 474065 15976 521455
rect 16040 498370 16068 587143
rect 16132 498438 16160 587182
rect 16212 586628 16264 586634
rect 16212 586570 16264 586576
rect 16224 499574 16252 586570
rect 16316 508337 16344 589222
rect 17132 587512 17184 587518
rect 17132 587454 17184 587460
rect 16396 587104 16448 587110
rect 16396 587046 16448 587052
rect 16302 508328 16358 508337
rect 16302 508263 16358 508272
rect 16224 499546 16344 499574
rect 16120 498432 16172 498438
rect 16120 498374 16172 498380
rect 16028 498364 16080 498370
rect 16028 498306 16080 498312
rect 16028 497616 16080 497622
rect 16028 497558 16080 497564
rect 15934 474056 15990 474065
rect 15934 473991 15990 474000
rect 15948 138310 15976 473991
rect 15936 138304 15988 138310
rect 15936 138246 15988 138252
rect 16040 106146 16068 497558
rect 16132 107438 16160 498374
rect 16316 498234 16344 499546
rect 16304 498228 16356 498234
rect 16304 498170 16356 498176
rect 16120 107432 16172 107438
rect 16120 107374 16172 107380
rect 16212 107024 16264 107030
rect 16212 106966 16264 106972
rect 16028 106140 16080 106146
rect 16028 106082 16080 106088
rect 15844 105664 15896 105670
rect 15844 105606 15896 105612
rect 16224 17678 16252 106966
rect 16316 105602 16344 498170
rect 16408 498098 16436 587046
rect 16488 586832 16540 586838
rect 16488 586774 16540 586780
rect 16396 498092 16448 498098
rect 16396 498034 16448 498040
rect 16500 496806 16528 586774
rect 17040 584792 17092 584798
rect 17040 584734 17092 584740
rect 16946 533760 17002 533769
rect 16946 533695 17002 533704
rect 16764 528624 16816 528630
rect 16764 528566 16816 528572
rect 16672 523796 16724 523802
rect 16672 523738 16724 523744
rect 16488 496800 16540 496806
rect 16488 496742 16540 496748
rect 16684 467158 16712 523738
rect 16672 467152 16724 467158
rect 16672 467094 16724 467100
rect 16684 140049 16712 467094
rect 16776 146985 16804 528566
rect 16856 523728 16908 523734
rect 16856 523670 16908 523676
rect 16868 468518 16896 523670
rect 16960 494834 16988 533695
rect 17052 498914 17080 584734
rect 17144 499050 17172 587454
rect 17236 532817 17264 622775
rect 17406 619984 17462 619993
rect 17406 619919 17462 619928
rect 17314 599992 17370 600001
rect 17314 599927 17370 599936
rect 17222 532808 17278 532817
rect 17222 532743 17278 532752
rect 17328 510610 17356 599927
rect 17420 531282 17448 619919
rect 17498 618216 17554 618225
rect 17498 618151 17554 618160
rect 17408 531276 17460 531282
rect 17408 531218 17460 531224
rect 17512 528193 17540 618151
rect 17604 536897 17632 626855
rect 17682 625968 17738 625977
rect 17682 625903 17738 625912
rect 17590 536888 17646 536897
rect 17590 536823 17646 536832
rect 17696 535945 17724 625903
rect 17866 623792 17922 623801
rect 17866 623727 17922 623736
rect 17774 621072 17830 621081
rect 17774 621007 17830 621016
rect 17682 535936 17738 535945
rect 17682 535871 17738 535880
rect 17590 532808 17646 532817
rect 17590 532743 17646 532752
rect 17498 528184 17554 528193
rect 17498 528119 17554 528128
rect 17512 527241 17540 528119
rect 17498 527232 17554 527241
rect 17498 527167 17554 527176
rect 17316 510604 17368 510610
rect 17316 510546 17368 510552
rect 17132 499044 17184 499050
rect 17132 498986 17184 498992
rect 17040 498908 17092 498914
rect 17040 498850 17092 498856
rect 16948 494828 17000 494834
rect 16948 494770 17000 494776
rect 16856 468512 16908 468518
rect 16856 468454 16908 468460
rect 16762 146976 16818 146985
rect 16762 146911 16818 146920
rect 16868 140865 16896 468454
rect 16960 144809 16988 494770
rect 17604 469878 17632 532743
rect 17696 472666 17724 535871
rect 17788 531049 17816 621007
rect 17880 533769 17908 623727
rect 19246 598360 19302 598369
rect 19246 598295 19302 598304
rect 19260 589286 19288 598295
rect 19248 589280 19300 589286
rect 19248 589222 19300 589228
rect 19154 587752 19210 587761
rect 19154 587687 19210 587696
rect 18604 587648 18656 587654
rect 18604 587590 18656 587596
rect 18420 587376 18472 587382
rect 18420 587318 18472 587324
rect 17866 533760 17922 533769
rect 17866 533695 17922 533704
rect 17774 531040 17830 531049
rect 17774 530975 17830 530984
rect 17788 523734 17816 530975
rect 17776 523728 17828 523734
rect 17776 523670 17828 523676
rect 17960 499656 18012 499662
rect 17960 499598 18012 499604
rect 17972 499526 18000 499598
rect 17960 499520 18012 499526
rect 17960 499462 18012 499468
rect 18328 498364 18380 498370
rect 18328 498306 18380 498312
rect 17684 472660 17736 472666
rect 17684 472602 17736 472608
rect 17592 469872 17644 469878
rect 17592 469814 17644 469820
rect 17132 195492 17184 195498
rect 17132 195434 17184 195440
rect 16946 144800 17002 144809
rect 16946 144735 17002 144744
rect 16854 140856 16910 140865
rect 16854 140791 16910 140800
rect 16670 140040 16726 140049
rect 16670 139975 16726 139984
rect 17038 120048 17094 120057
rect 17038 119983 17094 119992
rect 16488 107772 16540 107778
rect 16488 107714 16540 107720
rect 16396 106140 16448 106146
rect 16396 106082 16448 106088
rect 16304 105596 16356 105602
rect 16304 105538 16356 105544
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16408 17610 16436 106082
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 16500 16930 16528 107714
rect 17052 104854 17080 119983
rect 17144 107098 17172 195434
rect 17314 146976 17370 146985
rect 17314 146911 17370 146920
rect 17222 118416 17278 118425
rect 17222 118351 17278 118360
rect 17132 107092 17184 107098
rect 17132 107034 17184 107040
rect 17040 104848 17092 104854
rect 17040 104790 17092 104796
rect 17052 30025 17080 104790
rect 17038 30016 17094 30025
rect 17038 29951 17094 29960
rect 17144 19446 17172 107034
rect 17236 106282 17264 118351
rect 17224 106276 17276 106282
rect 17224 106218 17276 106224
rect 17236 28393 17264 106218
rect 17328 56953 17356 146911
rect 17406 146024 17462 146033
rect 17406 145959 17462 145968
rect 17314 56944 17370 56953
rect 17314 56879 17370 56888
rect 17420 56001 17448 145959
rect 17604 142905 17632 469814
rect 17696 146033 17724 472602
rect 17682 146024 17738 146033
rect 17682 145959 17738 145968
rect 17682 144800 17738 144809
rect 17682 144735 17738 144744
rect 17696 143857 17724 144735
rect 17682 143848 17738 143857
rect 17682 143783 17738 143792
rect 17590 142896 17646 142905
rect 17590 142831 17646 142840
rect 17604 142154 17632 142831
rect 17512 142126 17632 142154
rect 17406 55992 17462 56001
rect 17406 55927 17462 55936
rect 17512 52873 17540 142126
rect 17590 140040 17646 140049
rect 17590 139975 17646 139984
rect 17498 52864 17554 52873
rect 17498 52799 17554 52808
rect 17604 50017 17632 139975
rect 17696 53825 17724 143783
rect 17774 140856 17830 140865
rect 17774 140791 17830 140800
rect 17682 53816 17738 53825
rect 17682 53751 17738 53760
rect 17788 51105 17816 140791
rect 17868 138304 17920 138310
rect 17866 138272 17868 138281
rect 17920 138272 17922 138281
rect 17866 138207 17922 138216
rect 17774 51096 17830 51105
rect 17774 51031 17830 51040
rect 17590 50008 17646 50017
rect 17590 49943 17646 49952
rect 17880 48249 17908 138207
rect 18340 107930 18368 498306
rect 18432 497962 18460 587318
rect 18616 499526 18644 587590
rect 19064 584656 19116 584662
rect 19064 584598 19116 584604
rect 18788 531276 18840 531282
rect 18788 531218 18840 531224
rect 18800 529961 18828 531218
rect 18786 529952 18842 529961
rect 18786 529887 18842 529896
rect 18800 523802 18828 529887
rect 18788 523796 18840 523802
rect 18788 523738 18840 523744
rect 18604 499520 18656 499526
rect 18604 499462 18656 499468
rect 18616 499118 18644 499462
rect 18604 499112 18656 499118
rect 18604 499054 18656 499060
rect 19076 498166 19104 584598
rect 19064 498160 19116 498166
rect 19064 498102 19116 498108
rect 18420 497956 18472 497962
rect 18420 497898 18472 497904
rect 19168 497758 19196 587687
rect 19260 586498 19288 589222
rect 36634 587888 36690 587897
rect 36634 587823 36690 587832
rect 39578 587888 39634 587897
rect 39578 587823 39634 587832
rect 42798 587888 42854 587897
rect 42798 587823 42854 587832
rect 44178 587888 44234 587897
rect 44178 587823 44234 587832
rect 45282 587888 45338 587897
rect 45282 587823 45338 587832
rect 46846 587888 46902 587897
rect 46846 587823 46902 587832
rect 48134 587888 48190 587897
rect 48134 587823 48190 587832
rect 48686 587888 48742 587897
rect 48686 587823 48742 587832
rect 49790 587888 49846 587897
rect 49790 587823 49846 587832
rect 51078 587888 51134 587897
rect 51078 587823 51080 587832
rect 19800 587308 19852 587314
rect 19800 587250 19852 587256
rect 19708 586968 19760 586974
rect 19708 586910 19760 586916
rect 19248 586492 19300 586498
rect 19248 586434 19300 586440
rect 19338 536888 19394 536897
rect 19338 536823 19394 536832
rect 19352 528630 19380 536823
rect 19340 528624 19392 528630
rect 19340 528566 19392 528572
rect 19248 510604 19300 510610
rect 19248 510546 19300 510552
rect 19260 509969 19288 510546
rect 19246 509960 19302 509969
rect 19246 509895 19302 509904
rect 19260 498846 19288 509895
rect 19248 498840 19300 498846
rect 19248 498782 19300 498788
rect 19156 497752 19208 497758
rect 19156 497694 19208 497700
rect 19154 491192 19210 491201
rect 19154 491127 19210 491136
rect 19064 466472 19116 466478
rect 19064 466414 19116 466420
rect 18972 465112 19024 465118
rect 18972 465054 19024 465060
rect 18880 463752 18932 463758
rect 18880 463694 18932 463700
rect 18786 452840 18842 452849
rect 18786 452775 18842 452784
rect 18602 449848 18658 449857
rect 18602 449783 18658 449792
rect 18420 195560 18472 195566
rect 18420 195502 18472 195508
rect 18432 108118 18460 195502
rect 18512 195288 18564 195294
rect 18512 195230 18564 195236
rect 18420 108112 18472 108118
rect 18420 108054 18472 108060
rect 18340 107902 18460 107930
rect 18432 107273 18460 107902
rect 18524 107506 18552 195230
rect 18616 189038 18644 449783
rect 18696 195424 18748 195430
rect 18696 195366 18748 195372
rect 18604 189032 18656 189038
rect 18604 188974 18656 188980
rect 18708 107642 18736 195366
rect 18800 118153 18828 452775
rect 18786 118144 18842 118153
rect 18786 118079 18842 118088
rect 18696 107636 18748 107642
rect 18696 107578 18748 107584
rect 18512 107500 18564 107506
rect 18512 107442 18564 107448
rect 18788 107432 18840 107438
rect 18788 107374 18840 107380
rect 18418 107264 18474 107273
rect 18418 107199 18474 107208
rect 18328 106480 18380 106486
rect 18328 106422 18380 106428
rect 17866 48240 17922 48249
rect 17866 48175 17922 48184
rect 17222 28384 17278 28393
rect 17222 28319 17278 28328
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 18340 17338 18368 106422
rect 18432 18834 18460 107199
rect 18800 106486 18828 107374
rect 18892 107302 18920 463694
rect 18984 107438 19012 465054
rect 19076 107574 19104 466414
rect 19064 107568 19116 107574
rect 19064 107510 19116 107516
rect 18972 107432 19024 107438
rect 18972 107374 19024 107380
rect 18880 107296 18932 107302
rect 18880 107238 18932 107244
rect 18788 106480 18840 106486
rect 18788 106422 18840 106428
rect 18604 105732 18656 105738
rect 18604 105674 18656 105680
rect 18512 105664 18564 105670
rect 18512 105606 18564 105612
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18524 17814 18552 105606
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 18616 17746 18644 105674
rect 18696 105596 18748 105602
rect 18696 105538 18748 105544
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18708 17377 18736 105538
rect 18694 17368 18750 17377
rect 18328 17332 18380 17338
rect 18694 17303 18750 17312
rect 18328 17274 18380 17280
rect 18892 17134 18920 107238
rect 18984 17241 19012 107374
rect 19076 17950 19104 107510
rect 19168 107370 19196 491127
rect 19352 476814 19380 528566
rect 19430 508090 19486 508099
rect 19430 508025 19486 508034
rect 19444 478242 19472 508025
rect 19720 500002 19748 586910
rect 19708 499996 19760 500002
rect 19708 499938 19760 499944
rect 19720 499594 19748 499938
rect 19708 499588 19760 499594
rect 19708 499530 19760 499536
rect 19812 497554 19840 587250
rect 19984 587172 20036 587178
rect 19984 587114 20036 587120
rect 19892 586560 19944 586566
rect 19892 586502 19944 586508
rect 19904 497826 19932 586502
rect 19996 498030 20024 587114
rect 36648 586566 36676 587823
rect 39592 587382 39620 587823
rect 42812 587586 42840 587823
rect 44192 587790 44220 587823
rect 44180 587784 44232 587790
rect 44180 587726 44232 587732
rect 42800 587580 42852 587586
rect 42800 587522 42852 587528
rect 39580 587376 39632 587382
rect 39580 587318 39632 587324
rect 42812 587314 42840 587522
rect 42800 587308 42852 587314
rect 42800 587250 42852 587256
rect 44192 587042 44220 587726
rect 45296 587246 45324 587823
rect 46860 587382 46888 587823
rect 48148 587450 48176 587823
rect 48594 587752 48650 587761
rect 48594 587687 48650 587696
rect 48136 587444 48188 587450
rect 48136 587386 48188 587392
rect 46848 587376 46900 587382
rect 46848 587318 46900 587324
rect 45284 587240 45336 587246
rect 45284 587182 45336 587188
rect 46860 587110 46888 587318
rect 46848 587104 46900 587110
rect 46848 587046 46900 587052
rect 44180 587036 44232 587042
rect 44180 586978 44232 586984
rect 48148 586906 48176 587386
rect 48608 587178 48636 587687
rect 48596 587172 48648 587178
rect 48596 587114 48648 587120
rect 48136 586900 48188 586906
rect 48136 586842 48188 586848
rect 36636 586560 36688 586566
rect 36636 586502 36688 586508
rect 48700 584458 48728 587823
rect 49804 584526 49832 587823
rect 51132 587823 51134 587832
rect 52366 587888 52422 587897
rect 52366 587823 52422 587832
rect 53654 587888 53710 587897
rect 53654 587823 53710 587832
rect 53838 587888 53894 587897
rect 53838 587823 53894 587832
rect 55678 587888 55734 587897
rect 55678 587823 55734 587832
rect 56230 587888 56286 587897
rect 56230 587823 56286 587832
rect 59266 587888 59322 587897
rect 59266 587823 59322 587832
rect 60554 587888 60610 587897
rect 60554 587823 60610 587832
rect 61290 587888 61346 587897
rect 61290 587823 61346 587832
rect 62762 587888 62818 587897
rect 62762 587823 62818 587832
rect 63866 587888 63922 587897
rect 63866 587823 63922 587832
rect 64970 587888 65026 587897
rect 64970 587823 65026 587832
rect 66258 587888 66314 587897
rect 66258 587823 66314 587832
rect 67638 587888 67694 587897
rect 67638 587823 67694 587832
rect 68650 587888 68706 587897
rect 68650 587823 68706 587832
rect 69754 587888 69810 587897
rect 69754 587823 69756 587832
rect 51080 587794 51132 587800
rect 50066 587752 50122 587761
rect 50066 587687 50068 587696
rect 50120 587687 50122 587696
rect 50068 587658 50120 587664
rect 50080 586838 50108 587658
rect 51092 586974 51120 587794
rect 51080 586968 51132 586974
rect 51080 586910 51132 586916
rect 52380 586838 52408 587823
rect 52642 587752 52698 587761
rect 52642 587687 52698 587696
rect 50068 586832 50120 586838
rect 50068 586774 50120 586780
rect 51080 586832 51132 586838
rect 51080 586774 51132 586780
rect 52368 586832 52420 586838
rect 52368 586774 52420 586780
rect 51092 584662 51120 586774
rect 52656 586770 52684 587687
rect 52644 586764 52696 586770
rect 52644 586706 52696 586712
rect 51080 584656 51132 584662
rect 51080 584598 51132 584604
rect 52656 584594 52684 586706
rect 53668 584594 53696 587823
rect 53852 587654 53880 587823
rect 55692 587654 55720 587823
rect 53840 587648 53892 587654
rect 53840 587590 53892 587596
rect 55680 587648 55732 587654
rect 55680 587590 55732 587596
rect 53852 587246 53880 587590
rect 53840 587240 53892 587246
rect 53840 587182 53892 587188
rect 55692 586702 55720 587590
rect 55680 586696 55732 586702
rect 55680 586638 55732 586644
rect 56244 584662 56272 587823
rect 57058 587480 57114 587489
rect 57058 587415 57114 587424
rect 57072 586634 57100 587415
rect 57060 586628 57112 586634
rect 57060 586570 57112 586576
rect 59280 584730 59308 587823
rect 59818 587752 59874 587761
rect 59818 587687 59874 587696
rect 59832 586566 59860 587687
rect 60568 587518 60596 587823
rect 61304 587586 61332 587823
rect 62776 587790 62804 587823
rect 62764 587784 62816 587790
rect 62764 587726 62816 587732
rect 61292 587580 61344 587586
rect 61292 587522 61344 587528
rect 60556 587512 60608 587518
rect 60556 587454 60608 587460
rect 61842 587344 61898 587353
rect 63880 587314 63908 587823
rect 64984 587382 65012 587823
rect 65522 587752 65578 587761
rect 65522 587687 65578 587696
rect 65536 587489 65564 587687
rect 65522 587480 65578 587489
rect 65522 587415 65578 587424
rect 65982 587480 66038 587489
rect 66272 587450 66300 587823
rect 65982 587415 66038 587424
rect 66260 587444 66312 587450
rect 64972 587376 65024 587382
rect 63958 587344 64014 587353
rect 61842 587279 61898 587288
rect 63868 587308 63920 587314
rect 59820 586560 59872 586566
rect 59820 586502 59872 586508
rect 59832 584798 59860 586502
rect 61856 584798 61884 587279
rect 64972 587318 65024 587324
rect 63958 587279 64014 587288
rect 63868 587250 63920 587256
rect 63972 584866 64000 587279
rect 65996 584934 66024 587415
rect 66260 587386 66312 587392
rect 67652 587178 67680 587823
rect 68664 587722 68692 587823
rect 69808 587823 69810 587832
rect 71134 587888 71190 587897
rect 71134 587823 71190 587832
rect 72146 587888 72202 587897
rect 72146 587823 72202 587832
rect 73250 587888 73306 587897
rect 73250 587823 73306 587832
rect 73710 587888 73766 587897
rect 73710 587823 73766 587832
rect 74354 587888 74410 587897
rect 74354 587823 74410 587832
rect 76102 587888 76158 587897
rect 76102 587823 76158 587832
rect 77390 587888 77446 587897
rect 77390 587823 77446 587832
rect 78494 587888 78550 587897
rect 78494 587823 78550 587832
rect 79138 587888 79194 587897
rect 79138 587823 79194 587832
rect 81070 587888 81126 587897
rect 81070 587823 81126 587832
rect 83646 587888 83702 587897
rect 83646 587823 83702 587832
rect 88246 587888 88302 587897
rect 88246 587823 88302 587832
rect 91006 587888 91062 587897
rect 91006 587823 91062 587832
rect 93582 587888 93638 587897
rect 93582 587823 93638 587832
rect 96066 587888 96122 587897
rect 96066 587823 96122 587832
rect 98550 587888 98606 587897
rect 98550 587823 98606 587832
rect 100942 587888 100998 587897
rect 100942 587823 100998 587832
rect 103610 587888 103666 587897
rect 103610 587823 103666 587832
rect 105542 587888 105598 587897
rect 105542 587823 105598 587832
rect 108394 587888 108450 587897
rect 108394 587823 108450 587832
rect 111246 587888 111302 587897
rect 111246 587823 111302 587832
rect 113822 587888 113878 587897
rect 113822 587823 113878 587832
rect 114558 587888 114614 587897
rect 114558 587823 114614 587832
rect 118146 587888 118202 587897
rect 118146 587823 118202 587832
rect 120538 587888 120594 587897
rect 120538 587823 120594 587832
rect 125966 587888 126022 587897
rect 125966 587823 126022 587832
rect 69756 587794 69808 587800
rect 68652 587716 68704 587722
rect 68652 587658 68704 587664
rect 68558 587480 68614 587489
rect 68558 587415 68614 587424
rect 67640 587172 67692 587178
rect 67640 587114 67692 587120
rect 68572 585002 68600 587415
rect 71148 586838 71176 587823
rect 71136 586832 71188 586838
rect 71136 586774 71188 586780
rect 72160 586770 72188 587823
rect 73264 587246 73292 587823
rect 73252 587240 73304 587246
rect 73252 587182 73304 587188
rect 73724 586770 73752 587823
rect 74368 587654 74396 587823
rect 74356 587648 74408 587654
rect 74356 587590 74408 587596
rect 72148 586764 72200 586770
rect 72148 586706 72200 586712
rect 73712 586764 73764 586770
rect 73712 586706 73764 586712
rect 76116 586634 76144 587823
rect 76104 586628 76156 586634
rect 76104 586570 76156 586576
rect 77404 586566 77432 587823
rect 78508 586702 78536 587823
rect 79152 587518 79180 587823
rect 79140 587512 79192 587518
rect 79140 587454 79192 587460
rect 78496 586696 78548 586702
rect 78496 586638 78548 586644
rect 81084 586566 81112 587823
rect 83660 586906 83688 587823
rect 88260 586974 88288 587823
rect 88248 586968 88300 586974
rect 88248 586910 88300 586916
rect 83648 586900 83700 586906
rect 83648 586842 83700 586848
rect 91020 586838 91048 587823
rect 93596 587042 93624 587823
rect 96080 587110 96108 587823
rect 98564 587178 98592 587823
rect 100956 587246 100984 587823
rect 103624 587314 103652 587823
rect 103612 587308 103664 587314
rect 103612 587250 103664 587256
rect 100944 587240 100996 587246
rect 100944 587182 100996 587188
rect 98552 587172 98604 587178
rect 98552 587114 98604 587120
rect 96068 587104 96120 587110
rect 96068 587046 96120 587052
rect 93584 587036 93636 587042
rect 93584 586978 93636 586984
rect 91008 586832 91060 586838
rect 91008 586774 91060 586780
rect 77392 586560 77444 586566
rect 77392 586502 77444 586508
rect 81072 586560 81124 586566
rect 81072 586502 81124 586508
rect 105556 585070 105584 587823
rect 108408 585138 108436 587823
rect 111260 587382 111288 587823
rect 111248 587376 111300 587382
rect 111248 587318 111300 587324
rect 108396 585132 108448 585138
rect 108396 585074 108448 585080
rect 105544 585064 105596 585070
rect 105544 585006 105596 585012
rect 68560 584996 68612 585002
rect 68560 584938 68612 584944
rect 65984 584928 66036 584934
rect 65984 584870 66036 584876
rect 63960 584860 64012 584866
rect 63960 584802 64012 584808
rect 59820 584792 59872 584798
rect 59820 584734 59872 584740
rect 61844 584792 61896 584798
rect 61844 584734 61896 584740
rect 59268 584724 59320 584730
rect 59268 584666 59320 584672
rect 56232 584656 56284 584662
rect 56232 584598 56284 584604
rect 52644 584588 52696 584594
rect 52644 584530 52696 584536
rect 53656 584588 53708 584594
rect 53656 584530 53708 584536
rect 49792 584520 49844 584526
rect 49792 584462 49844 584468
rect 48688 584452 48740 584458
rect 48688 584394 48740 584400
rect 113836 584390 113864 587823
rect 113824 584384 113876 584390
rect 113824 584326 113876 584332
rect 114572 584322 114600 587823
rect 118160 584361 118188 587823
rect 120552 584497 120580 587823
rect 125980 587450 126008 587823
rect 125968 587444 126020 587450
rect 125968 587386 126020 587392
rect 156696 587444 156748 587450
rect 156696 587386 156748 587392
rect 156604 587308 156656 587314
rect 156604 587250 156656 587256
rect 122930 587072 122986 587081
rect 122930 587007 122986 587016
rect 122944 584633 122972 587007
rect 150716 586492 150768 586498
rect 150716 586434 150768 586440
rect 150728 585313 150756 586434
rect 150714 585304 150770 585313
rect 150714 585239 150770 585248
rect 122930 584624 122986 584633
rect 122930 584559 122986 584568
rect 120538 584488 120594 584497
rect 120538 584423 120594 584432
rect 118146 584352 118202 584361
rect 114560 584316 114612 584322
rect 118146 584287 118202 584296
rect 114560 584258 114612 584264
rect 20628 499996 20680 500002
rect 20628 499938 20680 499944
rect 20640 499186 20668 499938
rect 45374 499624 45430 499633
rect 45374 499559 45430 499568
rect 20628 499180 20680 499186
rect 20628 499122 20680 499128
rect 34520 498500 34572 498506
rect 34520 498442 34572 498448
rect 19984 498024 20036 498030
rect 19984 497966 20036 497972
rect 19892 497820 19944 497826
rect 19892 497762 19944 497768
rect 19996 497622 20024 497966
rect 34532 497894 34560 498442
rect 45388 498438 45416 499559
rect 51448 499180 51500 499186
rect 51448 499122 51500 499128
rect 44824 498432 44876 498438
rect 44824 498374 44876 498380
rect 45376 498432 45428 498438
rect 45376 498374 45428 498380
rect 37278 498128 37334 498137
rect 37278 498063 37334 498072
rect 41878 498128 41934 498137
rect 41878 498063 41934 498072
rect 43442 498128 43498 498137
rect 43442 498063 43498 498072
rect 34520 497888 34572 497894
rect 34520 497830 34572 497836
rect 36174 497856 36230 497865
rect 36174 497791 36230 497800
rect 37186 497856 37242 497865
rect 37186 497791 37188 497800
rect 36188 497758 36216 497791
rect 37240 497791 37242 497800
rect 37188 497762 37240 497768
rect 36176 497752 36228 497758
rect 36176 497694 36228 497700
rect 19984 497616 20036 497622
rect 22100 497616 22152 497622
rect 19984 497558 20036 497564
rect 22098 497584 22100 497593
rect 22152 497584 22154 497593
rect 19800 497548 19852 497554
rect 22098 497519 22154 497528
rect 19800 497490 19852 497496
rect 19812 496890 19840 497490
rect 20628 497208 20680 497214
rect 20628 497150 20680 497156
rect 19812 496862 19932 496890
rect 19800 496732 19852 496738
rect 19800 496674 19852 496680
rect 19432 478236 19484 478242
rect 19432 478178 19484 478184
rect 19340 476808 19392 476814
rect 19340 476750 19392 476756
rect 19708 451512 19760 451518
rect 19708 451454 19760 451460
rect 19616 195356 19668 195362
rect 19616 195298 19668 195304
rect 19248 108112 19300 108118
rect 19248 108054 19300 108060
rect 19260 107846 19288 108054
rect 19524 108044 19576 108050
rect 19524 107986 19576 107992
rect 19248 107840 19300 107846
rect 19248 107782 19300 107788
rect 19156 107364 19208 107370
rect 19156 107306 19208 107312
rect 19064 17944 19116 17950
rect 19064 17886 19116 17892
rect 19168 17513 19196 107306
rect 19154 17504 19210 17513
rect 19260 17474 19288 107782
rect 19432 107636 19484 107642
rect 19432 107578 19484 107584
rect 19444 106418 19472 107578
rect 19536 107166 19564 107986
rect 19628 107778 19656 195298
rect 19720 111790 19748 451454
rect 19708 111784 19760 111790
rect 19708 111726 19760 111732
rect 19812 108050 19840 496674
rect 19800 108044 19852 108050
rect 19800 107986 19852 107992
rect 19904 107930 19932 496862
rect 20640 496738 20668 497150
rect 34520 496800 34572 496806
rect 34520 496742 34572 496748
rect 20628 496732 20680 496738
rect 20628 496674 20680 496680
rect 19984 451444 20036 451450
rect 19984 451386 20036 451392
rect 19720 107902 19932 107930
rect 19616 107772 19668 107778
rect 19616 107714 19668 107720
rect 19616 107500 19668 107506
rect 19616 107442 19668 107448
rect 19524 107160 19576 107166
rect 19524 107102 19576 107108
rect 19432 106412 19484 106418
rect 19432 106354 19484 106360
rect 19154 17439 19210 17448
rect 19248 17468 19300 17474
rect 19248 17410 19300 17416
rect 19444 17406 19472 106354
rect 19432 17400 19484 17406
rect 19432 17342 19484 17348
rect 19536 17270 19564 107102
rect 19628 106350 19656 107442
rect 19720 107234 19748 107902
rect 19798 107536 19854 107545
rect 19798 107471 19854 107480
rect 19708 107228 19760 107234
rect 19708 107170 19760 107176
rect 19616 106344 19668 106350
rect 19616 106286 19668 106292
rect 19628 17882 19656 106286
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19524 17264 19576 17270
rect 18970 17232 19026 17241
rect 19524 17206 19576 17212
rect 19720 17202 19748 107170
rect 19812 106554 19840 107471
rect 19800 106548 19852 106554
rect 19800 106490 19852 106496
rect 19812 17649 19840 106490
rect 19996 33114 20024 451386
rect 34532 195566 34560 496742
rect 37292 491201 37320 498063
rect 39672 497956 39724 497962
rect 39672 497898 39724 497904
rect 38660 497752 38712 497758
rect 38660 497694 38712 497700
rect 37278 491192 37334 491201
rect 37278 491127 37334 491136
rect 37292 489258 37320 491127
rect 37280 489252 37332 489258
rect 37280 489194 37332 489200
rect 38672 465118 38700 497694
rect 39684 497049 39712 497898
rect 40592 497616 40644 497622
rect 40592 497558 40644 497564
rect 39670 497040 39726 497049
rect 39670 496975 39726 496984
rect 39684 496942 39712 496975
rect 39672 496936 39724 496942
rect 40604 496913 40632 497558
rect 39672 496878 39724 496884
rect 40590 496904 40646 496913
rect 40590 496839 40592 496848
rect 40644 496839 40646 496848
rect 40592 496810 40644 496816
rect 41892 494737 41920 498063
rect 42800 497820 42852 497826
rect 42800 497762 42852 497768
rect 41878 494728 41934 494737
rect 41878 494663 41934 494672
rect 41892 493474 41920 494663
rect 41880 493468 41932 493474
rect 41880 493410 41932 493416
rect 42812 466478 42840 497762
rect 43456 497554 43484 498063
rect 44178 497992 44234 498001
rect 44178 497927 44234 497936
rect 43444 497548 43496 497554
rect 43444 497490 43496 497496
rect 43456 497146 43484 497490
rect 44192 497214 44220 497927
rect 44836 497622 44864 498374
rect 51460 498137 51488 499122
rect 53840 499112 53892 499118
rect 53840 499054 53892 499060
rect 52184 498160 52236 498166
rect 46846 498128 46902 498137
rect 46846 498063 46848 498072
rect 46900 498063 46902 498072
rect 47582 498128 47638 498137
rect 47582 498063 47638 498072
rect 48686 498128 48742 498137
rect 48686 498063 48742 498072
rect 51446 498128 51502 498137
rect 51446 498063 51502 498072
rect 52182 498128 52184 498137
rect 53852 498137 53880 499054
rect 60740 499044 60792 499050
rect 60740 498986 60792 498992
rect 59544 498908 59596 498914
rect 59544 498850 59596 498856
rect 58164 498364 58216 498370
rect 58164 498306 58216 498312
rect 55864 498296 55916 498302
rect 55864 498238 55916 498244
rect 57888 498296 57940 498302
rect 57888 498238 57940 498244
rect 55876 498137 55904 498238
rect 57060 498228 57112 498234
rect 57060 498170 57112 498176
rect 52236 498128 52238 498137
rect 52182 498063 52238 498072
rect 53470 498128 53526 498137
rect 53470 498063 53526 498072
rect 53838 498128 53894 498137
rect 53838 498063 53894 498072
rect 55862 498128 55918 498137
rect 55862 498063 55918 498072
rect 46848 498034 46900 498040
rect 44824 497616 44876 497622
rect 44824 497558 44876 497564
rect 44180 497208 44232 497214
rect 44180 497150 44232 497156
rect 43444 497140 43496 497146
rect 43444 497082 43496 497088
rect 44180 496936 44232 496942
rect 44180 496878 44232 496884
rect 43444 496868 43496 496874
rect 43444 496810 43496 496816
rect 43456 474162 43484 496810
rect 43444 474156 43496 474162
rect 43444 474098 43496 474104
rect 42800 466472 42852 466478
rect 42800 466414 42852 466420
rect 43628 466472 43680 466478
rect 43628 466414 43680 466420
rect 43640 465798 43668 466414
rect 43628 465792 43680 465798
rect 43628 465734 43680 465740
rect 38660 465112 38712 465118
rect 38660 465054 38712 465060
rect 44192 463758 44220 496878
rect 46860 496874 46888 498034
rect 47596 497894 47624 498063
rect 48700 498030 48728 498063
rect 48688 498024 48740 498030
rect 48688 497966 48740 497972
rect 49608 498024 49660 498030
rect 49608 497966 49660 497972
rect 47584 497888 47636 497894
rect 47584 497830 47636 497836
rect 48228 497888 48280 497894
rect 48228 497830 48280 497836
rect 48240 496942 48268 497830
rect 49620 497554 49648 497966
rect 51460 497894 51488 498063
rect 51448 497888 51500 497894
rect 50250 497856 50306 497865
rect 51448 497830 51500 497836
rect 50250 497791 50306 497800
rect 49608 497548 49660 497554
rect 49608 497490 49660 497496
rect 50264 497078 50292 497791
rect 50252 497072 50304 497078
rect 50252 497014 50304 497020
rect 52196 497010 52224 498063
rect 53484 497962 53512 498063
rect 52460 497956 52512 497962
rect 52460 497898 52512 497904
rect 53472 497956 53524 497962
rect 53472 497898 53524 497904
rect 52472 497486 52500 497898
rect 53852 497758 53880 498063
rect 57072 497865 57100 498170
rect 57058 497856 57114 497865
rect 57900 497826 57928 498238
rect 58176 498001 58204 498306
rect 59556 498166 59584 498850
rect 59544 498160 59596 498166
rect 59542 498128 59544 498137
rect 59596 498128 59598 498137
rect 59542 498063 59598 498072
rect 60646 498128 60702 498137
rect 60752 498114 60780 498986
rect 78140 498166 78168 498197
rect 78128 498160 78180 498166
rect 60702 498086 60780 498114
rect 63682 498128 63738 498137
rect 60646 498063 60702 498072
rect 63682 498063 63738 498072
rect 64142 498128 64198 498137
rect 64142 498063 64198 498072
rect 67638 498128 67694 498137
rect 67638 498063 67694 498072
rect 71226 498128 71282 498137
rect 71226 498063 71282 498072
rect 71962 498128 72018 498137
rect 71962 498063 72018 498072
rect 73710 498128 73766 498137
rect 73710 498063 73766 498072
rect 73986 498128 74042 498137
rect 73986 498063 74042 498072
rect 78126 498128 78128 498137
rect 78180 498128 78182 498137
rect 78126 498063 78182 498072
rect 114466 498128 114522 498137
rect 114466 498063 114522 498072
rect 121366 498128 121422 498137
rect 121366 498063 121422 498072
rect 58162 497992 58218 498001
rect 58162 497927 58218 497936
rect 57058 497791 57114 497800
rect 57888 497820 57940 497826
rect 57888 497762 57940 497768
rect 53840 497752 53892 497758
rect 53840 497694 53892 497700
rect 60660 497690 60688 498063
rect 60648 497684 60700 497690
rect 60648 497626 60700 497632
rect 52460 497480 52512 497486
rect 52460 497422 52512 497428
rect 62764 497208 62816 497214
rect 62764 497150 62816 497156
rect 61844 497140 61896 497146
rect 61844 497082 61896 497088
rect 61856 497049 61884 497082
rect 61842 497040 61898 497049
rect 52184 497004 52236 497010
rect 52184 496946 52236 496952
rect 52460 497004 52512 497010
rect 61842 496975 61898 496984
rect 52460 496946 52512 496952
rect 48228 496936 48280 496942
rect 48228 496878 48280 496884
rect 48318 496904 48374 496913
rect 46848 496868 46900 496874
rect 48318 496839 48374 496848
rect 50986 496904 51042 496913
rect 50986 496839 51042 496848
rect 46848 496810 46900 496816
rect 48332 493542 48360 496839
rect 48320 493536 48372 493542
rect 48320 493478 48372 493484
rect 44180 463752 44232 463758
rect 44180 463694 44232 463700
rect 44640 463752 44692 463758
rect 44640 463694 44692 463700
rect 44652 463078 44680 463694
rect 44640 463072 44692 463078
rect 44640 463014 44692 463020
rect 51000 453558 51028 496839
rect 50988 453552 51040 453558
rect 50988 453494 51040 453500
rect 48964 451716 49016 451722
rect 48964 451658 49016 451664
rect 34520 195560 34572 195566
rect 34520 195502 34572 195508
rect 48976 193866 49004 451658
rect 52472 195498 52500 496946
rect 53746 496904 53802 496913
rect 53746 496839 53802 496848
rect 56506 496904 56562 496913
rect 56506 496839 56562 496848
rect 59266 496904 59322 496913
rect 59266 496839 59322 496848
rect 53760 471306 53788 496839
rect 53748 471300 53800 471306
rect 53748 471242 53800 471248
rect 56520 453490 56548 496839
rect 56508 453484 56560 453490
rect 56508 453426 56560 453432
rect 59280 453422 59308 496839
rect 61856 490754 61884 496975
rect 62776 496913 62804 497150
rect 62026 496904 62082 496913
rect 62026 496839 62082 496848
rect 62762 496904 62818 496913
rect 62762 496839 62818 496848
rect 61844 490748 61896 490754
rect 61844 490690 61896 490696
rect 59268 453416 59320 453422
rect 59268 453358 59320 453364
rect 62040 453354 62068 496839
rect 62776 487150 62804 496839
rect 63696 496126 63724 498063
rect 64156 497622 64184 498063
rect 64144 497616 64196 497622
rect 64144 497558 64196 497564
rect 63684 496120 63736 496126
rect 63684 496062 63736 496068
rect 64156 489870 64184 497558
rect 67652 497554 67680 498063
rect 69664 497888 69716 497894
rect 69664 497830 69716 497836
rect 67640 497548 67692 497554
rect 67640 497490 67692 497496
rect 68928 497548 68980 497554
rect 68928 497490 68980 497496
rect 68282 497176 68338 497185
rect 68282 497111 68338 497120
rect 68296 497078 68324 497111
rect 68284 497072 68336 497078
rect 66258 497040 66314 497049
rect 68284 497014 68336 497020
rect 66258 496975 66314 496984
rect 66272 496942 66300 496975
rect 66260 496936 66312 496942
rect 65522 496904 65578 496913
rect 65522 496839 65524 496848
rect 65576 496839 65578 496848
rect 66166 496904 66222 496913
rect 66260 496878 66312 496884
rect 66904 496936 66956 496942
rect 66904 496878 66956 496884
rect 66166 496839 66222 496848
rect 65524 496810 65576 496816
rect 64144 489864 64196 489870
rect 64144 489806 64196 489812
rect 62764 487144 62816 487150
rect 62764 487086 62816 487092
rect 65536 465594 65564 496810
rect 66180 481030 66208 496839
rect 66916 487898 66944 496878
rect 66904 487892 66956 487898
rect 66904 487834 66956 487840
rect 66168 481024 66220 481030
rect 66168 480966 66220 480972
rect 68296 476950 68324 497014
rect 68940 496942 68968 497490
rect 68928 496936 68980 496942
rect 68558 496904 68614 496913
rect 69676 496913 69704 497830
rect 71240 497486 71268 498063
rect 71976 497962 72004 498063
rect 71964 497956 72016 497962
rect 71964 497898 72016 497904
rect 70400 497480 70452 497486
rect 70400 497422 70452 497428
rect 71228 497480 71280 497486
rect 71228 497422 71280 497428
rect 70412 497010 70440 497422
rect 71976 497078 72004 497898
rect 73160 497752 73212 497758
rect 73158 497720 73160 497729
rect 73212 497720 73214 497729
rect 73158 497655 73214 497664
rect 71964 497072 72016 497078
rect 71964 497014 72016 497020
rect 70400 497004 70452 497010
rect 70400 496946 70452 496952
rect 68928 496878 68980 496884
rect 69662 496904 69718 496913
rect 68558 496839 68614 496848
rect 69662 496839 69718 496848
rect 71686 496904 71742 496913
rect 71686 496839 71742 496848
rect 68572 490686 68600 496839
rect 68560 490680 68612 490686
rect 68560 490622 68612 490628
rect 68284 476944 68336 476950
rect 68284 476886 68336 476892
rect 69676 470558 69704 496839
rect 71700 482458 71728 496839
rect 73724 492046 73752 498063
rect 74000 497826 74028 498063
rect 76562 497992 76618 498001
rect 76562 497927 76618 497936
rect 75182 497856 75238 497865
rect 73988 497820 74040 497826
rect 75182 497791 75238 497800
rect 73988 497762 74040 497768
rect 73802 496904 73858 496913
rect 73802 496839 73858 496848
rect 73712 492040 73764 492046
rect 73712 491982 73764 491988
rect 71688 482452 71740 482458
rect 71688 482394 71740 482400
rect 73816 475454 73844 496839
rect 74000 485790 74028 497762
rect 73988 485784 74040 485790
rect 73988 485726 74040 485732
rect 73804 475448 73856 475454
rect 73804 475390 73856 475396
rect 75196 471986 75224 497791
rect 76576 472734 76604 497927
rect 78140 497146 78168 498063
rect 79416 497684 79468 497690
rect 79416 497626 79468 497632
rect 78128 497140 78180 497146
rect 78128 497082 78180 497088
rect 79324 497140 79376 497146
rect 79324 497082 79376 497088
rect 76838 496904 76894 496913
rect 76838 496839 76894 496848
rect 78586 496904 78642 496913
rect 78586 496839 78642 496848
rect 76852 490618 76880 496839
rect 76840 490612 76892 490618
rect 76840 490554 76892 490560
rect 78600 489190 78628 496839
rect 78588 489184 78640 489190
rect 78588 489126 78640 489132
rect 76564 472728 76616 472734
rect 76564 472670 76616 472676
rect 75184 471980 75236 471986
rect 75184 471922 75236 471928
rect 69664 470552 69716 470558
rect 69664 470494 69716 470500
rect 65524 465588 65576 465594
rect 65524 465530 65576 465536
rect 66260 465588 66312 465594
rect 66260 465530 66312 465536
rect 66272 465118 66300 465530
rect 66260 465112 66312 465118
rect 66260 465054 66312 465060
rect 62028 453348 62080 453354
rect 62028 453290 62080 453296
rect 52460 195492 52512 195498
rect 52460 195434 52512 195440
rect 66272 195430 66300 465054
rect 79336 464982 79364 497082
rect 79428 496913 79456 497626
rect 106094 497176 106150 497185
rect 106094 497111 106150 497120
rect 79414 496904 79470 496913
rect 79414 496839 79470 496848
rect 81346 496904 81402 496913
rect 81346 496839 81402 496848
rect 84106 496904 84162 496913
rect 84106 496839 84162 496848
rect 86866 496904 86922 496913
rect 86866 496839 86922 496848
rect 88246 496904 88302 496913
rect 88246 496839 88302 496848
rect 91006 496904 91062 496913
rect 91006 496839 91062 496848
rect 93766 496904 93822 496913
rect 93766 496839 93822 496848
rect 96526 496904 96582 496913
rect 96526 496839 96582 496848
rect 99286 496904 99342 496913
rect 99286 496839 99342 496848
rect 100942 496904 100998 496913
rect 100942 496839 100998 496848
rect 104806 496904 104862 496913
rect 104806 496839 104862 496848
rect 79428 466478 79456 496839
rect 81360 480962 81388 496839
rect 84120 482390 84148 496839
rect 86880 483750 86908 496839
rect 88260 487830 88288 496839
rect 88248 487824 88300 487830
rect 88248 487766 88300 487772
rect 91020 486538 91048 496839
rect 91008 486532 91060 486538
rect 91008 486474 91060 486480
rect 86868 483744 86920 483750
rect 86868 483686 86920 483692
rect 84108 482384 84160 482390
rect 84108 482326 84160 482332
rect 81348 480956 81400 480962
rect 81348 480898 81400 480904
rect 93780 479534 93808 496839
rect 96540 485110 96568 496839
rect 96528 485104 96580 485110
rect 96528 485046 96580 485052
rect 93768 479528 93820 479534
rect 93768 479470 93820 479476
rect 99300 475386 99328 496839
rect 100956 493406 100984 496839
rect 100944 493400 100996 493406
rect 100944 493342 100996 493348
rect 104820 478310 104848 496839
rect 106108 494902 106136 497111
rect 108854 496904 108910 496913
rect 108854 496839 108910 496848
rect 111706 496904 111762 496913
rect 111706 496839 111762 496848
rect 106096 494896 106148 494902
rect 106096 494838 106148 494844
rect 108868 491978 108896 496839
rect 108856 491972 108908 491978
rect 108856 491914 108908 491920
rect 104808 478304 104860 478310
rect 104808 478246 104860 478252
rect 99288 475380 99340 475386
rect 99288 475322 99340 475328
rect 80704 474768 80756 474774
rect 80704 474710 80756 474716
rect 79416 466472 79468 466478
rect 79416 466414 79468 466420
rect 80060 466472 80112 466478
rect 80060 466414 80112 466420
rect 79324 464976 79376 464982
rect 79324 464918 79376 464924
rect 66260 195424 66312 195430
rect 66260 195366 66312 195372
rect 80072 195294 80100 466414
rect 80152 464976 80204 464982
rect 80152 464918 80204 464924
rect 80164 463758 80192 464918
rect 80152 463752 80204 463758
rect 80152 463694 80204 463700
rect 80164 195362 80192 463694
rect 80716 457842 80744 474710
rect 80704 457836 80756 457842
rect 80704 457778 80756 457784
rect 111720 454714 111748 496839
rect 114480 474094 114508 498063
rect 115846 496904 115902 496913
rect 115846 496839 115902 496848
rect 118606 496904 118662 496913
rect 118606 496839 118662 496848
rect 115860 476882 115888 496839
rect 115848 476876 115900 476882
rect 115848 476818 115900 476824
rect 114468 474088 114520 474094
rect 114468 474030 114520 474036
rect 118620 469946 118648 496839
rect 118608 469940 118660 469946
rect 118608 469882 118660 469888
rect 121380 463010 121408 498063
rect 124126 496904 124182 496913
rect 124126 496839 124182 496848
rect 126886 496904 126942 496913
rect 126886 496839 126942 496848
rect 124140 464370 124168 496839
rect 126900 465730 126928 496839
rect 126888 465724 126940 465730
rect 126888 465666 126940 465672
rect 124128 464364 124180 464370
rect 124128 464306 124180 464312
rect 121368 463004 121420 463010
rect 121368 462946 121420 462952
rect 156616 460290 156644 587250
rect 156708 465769 156736 587386
rect 156788 587240 156840 587246
rect 156788 587182 156840 587188
rect 156800 485246 156828 587182
rect 157352 586498 157380 674834
rect 158718 668672 158774 668681
rect 158718 668607 158774 668616
rect 158076 587172 158128 587178
rect 158076 587114 158128 587120
rect 157984 586764 158036 586770
rect 157984 586706 158036 586712
rect 157340 586492 157392 586498
rect 157340 586434 157392 586440
rect 157352 585721 157380 586434
rect 157338 585712 157394 585721
rect 157338 585647 157394 585656
rect 156788 485240 156840 485246
rect 156788 485182 156840 485188
rect 157996 467226 158024 586706
rect 158088 472802 158116 587114
rect 158168 587036 158220 587042
rect 158168 586978 158220 586984
rect 158180 486606 158208 586978
rect 158260 586900 158312 586906
rect 158260 586842 158312 586848
rect 158272 487966 158300 586842
rect 158732 579193 158760 668607
rect 162124 587376 162176 587382
rect 162124 587318 162176 587324
rect 159456 587104 159508 587110
rect 159456 587046 159508 587052
rect 159364 586968 159416 586974
rect 159364 586910 159416 586916
rect 158718 579184 158774 579193
rect 158718 579119 158774 579128
rect 158260 487960 158312 487966
rect 158260 487902 158312 487908
rect 158168 486600 158220 486606
rect 158168 486542 158220 486548
rect 158076 472796 158128 472802
rect 158076 472738 158128 472744
rect 157984 467220 158036 467226
rect 157984 467162 158036 467168
rect 156694 465760 156750 465769
rect 156694 465695 156750 465704
rect 156604 460284 156656 460290
rect 156604 460226 156656 460232
rect 157984 455048 158036 455054
rect 157984 454990 158036 454996
rect 111708 454708 111760 454714
rect 111708 454650 111760 454656
rect 156604 450900 156656 450906
rect 156604 450842 156656 450848
rect 150990 196072 151046 196081
rect 150990 196007 150992 196016
rect 151044 196007 151046 196016
rect 150992 195978 151044 195984
rect 80152 195356 80204 195362
rect 80152 195298 80204 195304
rect 80060 195288 80112 195294
rect 80060 195230 80112 195236
rect 48964 193860 49016 193866
rect 48964 193802 49016 193808
rect 50802 109576 50858 109585
rect 50802 109511 50858 109520
rect 56046 109576 56102 109585
rect 56046 109511 56102 109520
rect 61106 109576 61162 109585
rect 61106 109511 61162 109520
rect 106002 109576 106058 109585
rect 106002 109511 106058 109520
rect 108578 109576 108634 109585
rect 108578 109511 108634 109520
rect 48318 109032 48374 109041
rect 48318 108967 48374 108976
rect 48332 108322 48360 108967
rect 50816 108390 50844 109511
rect 53654 108760 53710 108769
rect 53654 108695 53710 108704
rect 53668 108458 53696 108695
rect 56060 108526 56088 109511
rect 61120 108594 61148 109511
rect 68374 109032 68430 109041
rect 68374 108967 68430 108976
rect 100942 109032 100998 109041
rect 100942 108967 100998 108976
rect 68388 108662 68416 108967
rect 100956 108730 100984 108967
rect 106016 108798 106044 109511
rect 108592 108866 108620 109511
rect 111062 109032 111118 109041
rect 111062 108967 111118 108976
rect 113454 109032 113510 109041
rect 113454 108967 113456 108976
rect 111076 108934 111104 108967
rect 113508 108967 113510 108976
rect 113456 108938 113508 108944
rect 111064 108928 111116 108934
rect 111064 108870 111116 108876
rect 108580 108860 108632 108866
rect 108580 108802 108632 108808
rect 106004 108792 106056 108798
rect 106004 108734 106056 108740
rect 100944 108724 100996 108730
rect 100944 108666 100996 108672
rect 68376 108656 68428 108662
rect 68376 108598 68428 108604
rect 61108 108588 61160 108594
rect 61108 108530 61160 108536
rect 56048 108520 56100 108526
rect 56048 108462 56100 108468
rect 53656 108452 53708 108458
rect 53656 108394 53708 108400
rect 50804 108384 50856 108390
rect 50804 108326 50856 108332
rect 48320 108316 48372 108322
rect 48320 108258 48372 108264
rect 50160 107704 50212 107710
rect 50160 107646 50212 107652
rect 50172 107574 50200 107646
rect 59636 107636 59688 107642
rect 59636 107578 59688 107584
rect 63592 107636 63644 107642
rect 63592 107578 63644 107584
rect 36912 107568 36964 107574
rect 35898 107536 35954 107545
rect 35898 107471 35954 107480
rect 36910 107536 36912 107545
rect 50160 107568 50212 107574
rect 36964 107536 36966 107545
rect 36910 107471 36966 107480
rect 38106 107536 38162 107545
rect 38106 107471 38162 107480
rect 39578 107536 39634 107545
rect 39578 107471 39634 107480
rect 40498 107536 40554 107545
rect 40498 107471 40554 107480
rect 43166 107536 43222 107545
rect 43166 107471 43168 107480
rect 35912 107438 35940 107471
rect 35900 107432 35952 107438
rect 35900 107374 35952 107380
rect 38120 107370 38148 107471
rect 38108 107364 38160 107370
rect 38108 107306 38160 107312
rect 39592 107302 39620 107471
rect 39580 107296 39632 107302
rect 39580 107238 39632 107244
rect 40512 106554 40540 107471
rect 43220 107471 43222 107480
rect 44270 107536 44326 107545
rect 44270 107471 44326 107480
rect 45374 107536 45430 107545
rect 45374 107471 45430 107480
rect 46570 107536 46626 107545
rect 46570 107471 46626 107480
rect 47582 107536 47638 107545
rect 47582 107471 47638 107480
rect 48778 107536 48834 107545
rect 48778 107471 48834 107480
rect 50158 107536 50160 107545
rect 59648 107545 59676 107578
rect 63604 107545 63632 107578
rect 68652 107568 68704 107574
rect 50212 107536 50214 107545
rect 50158 107471 50214 107480
rect 51262 107536 51318 107545
rect 51262 107471 51318 107480
rect 52366 107536 52422 107545
rect 52366 107471 52422 107480
rect 53470 107536 53526 107545
rect 53470 107471 53526 107480
rect 59634 107536 59690 107545
rect 59634 107471 59690 107480
rect 60554 107536 60610 107545
rect 60554 107471 60610 107480
rect 61658 107536 61714 107545
rect 62578 107536 62634 107545
rect 61658 107471 61660 107480
rect 43168 107442 43220 107448
rect 44284 107234 44312 107471
rect 45388 107370 45416 107471
rect 44364 107364 44416 107370
rect 44364 107306 44416 107312
rect 45376 107364 45428 107370
rect 45376 107306 45428 107312
rect 44272 107228 44324 107234
rect 44272 107170 44324 107176
rect 44180 107160 44232 107166
rect 44180 107102 44232 107108
rect 40500 106548 40552 106554
rect 40500 106490 40552 106496
rect 42800 106548 42852 106554
rect 42800 106490 42852 106496
rect 42812 106146 42840 106490
rect 44192 106214 44220 107102
rect 44284 106826 44312 107170
rect 44272 106820 44324 106826
rect 44272 106762 44324 106768
rect 44376 106486 44404 107306
rect 46584 107302 46612 107471
rect 46572 107296 46624 107302
rect 46572 107238 46624 107244
rect 44364 106480 44416 106486
rect 44364 106422 44416 106428
rect 46584 106418 46612 107238
rect 47596 107166 47624 107471
rect 48792 107234 48820 107471
rect 48780 107228 48832 107234
rect 48780 107170 48832 107176
rect 47584 107160 47636 107166
rect 47584 107102 47636 107108
rect 48792 106554 48820 107170
rect 51276 107030 51304 107471
rect 52276 107432 52328 107438
rect 52276 107374 52328 107380
rect 52288 107030 52316 107374
rect 52380 107098 52408 107471
rect 52368 107092 52420 107098
rect 52368 107034 52420 107040
rect 51264 107024 51316 107030
rect 51264 106966 51316 106972
rect 52276 107024 52328 107030
rect 52276 106966 52328 106972
rect 53484 106962 53512 107471
rect 55126 107128 55182 107137
rect 55770 107128 55826 107137
rect 55182 107086 55352 107114
rect 55126 107063 55182 107072
rect 53472 106956 53524 106962
rect 53472 106898 53524 106904
rect 48780 106548 48832 106554
rect 48780 106490 48832 106496
rect 55324 106418 55352 107086
rect 55770 107063 55826 107072
rect 59360 107092 59412 107098
rect 55784 106486 55812 107063
rect 59360 107034 59412 107040
rect 55772 106480 55824 106486
rect 55772 106422 55824 106428
rect 46572 106412 46624 106418
rect 46572 106354 46624 106360
rect 55312 106412 55364 106418
rect 55312 106354 55364 106360
rect 44180 106208 44232 106214
rect 44180 106150 44232 106156
rect 42800 106140 42852 106146
rect 42800 106082 42852 106088
rect 55324 105738 55352 106354
rect 55312 105732 55364 105738
rect 55312 105674 55364 105680
rect 55784 105670 55812 106422
rect 59372 106350 59400 107034
rect 59648 106894 59676 107471
rect 60568 107098 60596 107471
rect 61712 107471 61714 107480
rect 61752 107500 61804 107506
rect 61660 107442 61712 107448
rect 62578 107471 62634 107480
rect 63590 107536 63646 107545
rect 63590 107471 63646 107480
rect 63866 107536 63922 107545
rect 63866 107471 63922 107480
rect 65154 107536 65210 107545
rect 65154 107471 65210 107480
rect 66258 107536 66314 107545
rect 66258 107471 66314 107480
rect 67638 107536 67694 107545
rect 67638 107471 67694 107480
rect 68650 107536 68652 107545
rect 73712 107568 73764 107574
rect 68704 107536 68706 107545
rect 68650 107471 68706 107480
rect 69754 107536 69810 107545
rect 69754 107471 69810 107480
rect 71226 107536 71282 107545
rect 71226 107471 71282 107480
rect 72146 107536 72202 107545
rect 72146 107471 72202 107480
rect 73250 107536 73306 107545
rect 73250 107471 73306 107480
rect 73710 107536 73712 107545
rect 73764 107536 73766 107545
rect 73710 107471 73766 107480
rect 74354 107536 74410 107545
rect 74354 107471 74410 107480
rect 75642 107536 75698 107545
rect 75642 107471 75644 107480
rect 61752 107442 61804 107448
rect 61764 107409 61792 107442
rect 61750 107400 61806 107409
rect 61750 107335 61806 107344
rect 60556 107092 60608 107098
rect 60556 107034 60608 107040
rect 59636 106888 59688 106894
rect 59636 106830 59688 106836
rect 62592 106826 62620 107471
rect 63880 107370 63908 107471
rect 63868 107364 63920 107370
rect 63868 107306 63920 107312
rect 65168 107302 65196 107471
rect 65156 107296 65208 107302
rect 65156 107238 65208 107244
rect 66272 107166 66300 107471
rect 67652 107234 67680 107471
rect 69768 107438 69796 107471
rect 69756 107432 69808 107438
rect 69756 107374 69808 107380
rect 67640 107228 67692 107234
rect 67640 107170 67692 107176
rect 66260 107160 66312 107166
rect 66260 107102 66312 107108
rect 71240 107030 71268 107471
rect 71228 107024 71280 107030
rect 71228 106966 71280 106972
rect 72160 106962 72188 107471
rect 72148 106956 72200 106962
rect 72148 106898 72200 106904
rect 62580 106820 62632 106826
rect 62580 106762 62632 106768
rect 73264 106418 73292 107471
rect 74368 106486 74396 107471
rect 75696 107471 75698 107480
rect 76102 107536 76158 107545
rect 76102 107471 76104 107480
rect 75644 107442 75696 107448
rect 76156 107471 76158 107480
rect 77666 107536 77722 107545
rect 77666 107471 77722 107480
rect 78494 107536 78550 107545
rect 78494 107471 78550 107480
rect 79138 107536 79194 107545
rect 79138 107471 79194 107480
rect 86038 107536 86094 107545
rect 86038 107471 86094 107480
rect 88246 107536 88302 107545
rect 88246 107471 88302 107480
rect 93582 107536 93638 107545
rect 93582 107471 93638 107480
rect 98550 107536 98606 107545
rect 98550 107471 98606 107480
rect 120998 107536 121054 107545
rect 120998 107471 121054 107480
rect 123390 107536 123446 107545
rect 123390 107471 123446 107480
rect 76104 107442 76156 107448
rect 77680 106894 77708 107471
rect 78508 107438 78536 107471
rect 78496 107432 78548 107438
rect 78496 107374 78548 107380
rect 79152 107098 79180 107471
rect 86052 107370 86080 107471
rect 86040 107364 86092 107370
rect 86040 107306 86092 107312
rect 88260 107302 88288 107471
rect 88248 107296 88300 107302
rect 88248 107238 88300 107244
rect 93596 107234 93624 107471
rect 93584 107228 93636 107234
rect 93584 107170 93636 107176
rect 79140 107092 79192 107098
rect 79140 107034 79192 107040
rect 98564 107030 98592 107471
rect 121012 107166 121040 107471
rect 121000 107160 121052 107166
rect 121000 107102 121052 107108
rect 123404 107098 123432 107471
rect 156616 107302 156644 450842
rect 156696 450832 156748 450838
rect 156696 450774 156748 450780
rect 156604 107296 156656 107302
rect 156604 107238 156656 107244
rect 123392 107092 123444 107098
rect 123392 107034 123444 107040
rect 156708 107030 156736 450774
rect 157340 196036 157392 196042
rect 157340 195978 157392 195984
rect 98552 107024 98604 107030
rect 98552 106966 98604 106972
rect 156696 107024 156748 107030
rect 156696 106966 156748 106972
rect 77668 106888 77720 106894
rect 77668 106830 77720 106836
rect 74356 106480 74408 106486
rect 74356 106422 74408 106428
rect 73252 106412 73304 106418
rect 73252 106354 73304 106360
rect 59360 106344 59412 106350
rect 57058 106312 57114 106321
rect 59360 106286 59412 106292
rect 157352 106282 157380 195978
rect 57058 106247 57114 106256
rect 150808 106276 150860 106282
rect 55772 105664 55824 105670
rect 55772 105606 55824 105612
rect 57072 105602 57100 106247
rect 150808 106218 150860 106224
rect 157340 106276 157392 106282
rect 157340 106218 157392 106224
rect 57060 105596 57112 105602
rect 57060 105538 57112 105544
rect 150820 105369 150848 106218
rect 150806 105360 150862 105369
rect 150806 105295 150862 105304
rect 19984 33108 20036 33114
rect 19984 33050 20036 33056
rect 52366 19544 52422 19553
rect 52366 19479 52422 19488
rect 53470 19544 53526 19553
rect 53470 19479 53526 19488
rect 55954 19544 56010 19553
rect 55954 19479 56010 19488
rect 52380 19446 52408 19479
rect 52368 19440 52420 19446
rect 52368 19382 52420 19388
rect 50894 18728 50950 18737
rect 50894 18663 50950 18672
rect 50908 18630 50936 18663
rect 50896 18624 50948 18630
rect 50896 18566 50948 18572
rect 36544 17944 36596 17950
rect 36542 17912 36544 17921
rect 36596 17912 36598 17921
rect 36542 17847 36598 17856
rect 43074 17912 43130 17921
rect 43074 17847 43130 17856
rect 44178 17912 44234 17921
rect 44178 17847 44234 17856
rect 45374 17912 45430 17921
rect 45374 17847 45430 17856
rect 46662 17912 46718 17921
rect 46662 17847 46718 17856
rect 47582 17912 47638 17921
rect 47582 17847 47638 17856
rect 48686 17912 48742 17921
rect 48686 17847 48742 17856
rect 50158 17912 50214 17921
rect 50158 17847 50214 17856
rect 51446 17912 51502 17921
rect 51446 17847 51502 17856
rect 19798 17640 19854 17649
rect 19798 17575 19854 17584
rect 38658 17232 38714 17241
rect 18970 17167 19026 17176
rect 19708 17196 19760 17202
rect 38658 17167 38714 17176
rect 19708 17138 19760 17144
rect 38672 17134 38700 17167
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 38660 17128 38712 17134
rect 38660 17070 38712 17076
rect 43088 17066 43116 17847
rect 44192 17134 44220 17847
rect 45388 17202 45416 17847
rect 46676 17270 46704 17847
rect 47596 17542 47624 17847
rect 48700 17610 48728 17847
rect 48688 17604 48740 17610
rect 48688 17546 48740 17552
rect 49608 17604 49660 17610
rect 49608 17546 49660 17552
rect 47584 17536 47636 17542
rect 47584 17478 47636 17484
rect 48228 17536 48280 17542
rect 48228 17478 48280 17484
rect 48240 17338 48268 17478
rect 49620 17406 49648 17546
rect 50172 17542 50200 17847
rect 51460 17678 51488 17847
rect 51448 17672 51500 17678
rect 51448 17614 51500 17620
rect 50160 17536 50212 17542
rect 50160 17478 50212 17484
rect 49608 17400 49660 17406
rect 49608 17342 49660 17348
rect 48228 17332 48280 17338
rect 48228 17274 48280 17280
rect 46664 17264 46716 17270
rect 46664 17206 46716 17212
rect 45376 17196 45428 17202
rect 45376 17138 45428 17144
rect 44180 17128 44232 17134
rect 44180 17070 44232 17076
rect 43076 17060 43128 17066
rect 43076 17002 43128 17008
rect 51460 16998 51488 17614
rect 51448 16992 51500 16998
rect 51448 16934 51500 16940
rect 16488 16924 16540 16930
rect 16488 16866 16540 16872
rect 52380 16726 52408 19382
rect 53484 19378 53512 19479
rect 53472 19372 53524 19378
rect 53472 19314 53524 19320
rect 53484 17610 53512 19314
rect 53654 18728 53710 18737
rect 53654 18663 53656 18672
rect 53708 18663 53710 18672
rect 53656 18634 53708 18640
rect 55968 17814 55996 19479
rect 103704 19304 103756 19310
rect 95974 19272 96030 19281
rect 95974 19207 96030 19216
rect 100942 19272 100998 19281
rect 100942 19207 100944 19216
rect 95988 19174 96016 19207
rect 100996 19207 100998 19216
rect 103702 19272 103704 19281
rect 103756 19272 103758 19281
rect 103702 19207 103758 19216
rect 100944 19178 100996 19184
rect 95976 19168 96028 19174
rect 86038 19136 86094 19145
rect 86038 19071 86094 19080
rect 91006 19136 91062 19145
rect 95976 19110 96028 19116
rect 91006 19071 91008 19080
rect 86052 19038 86080 19071
rect 91060 19071 91062 19080
rect 91008 19042 91060 19048
rect 86040 19032 86092 19038
rect 76102 19000 76158 19009
rect 76102 18935 76158 18944
rect 81070 19000 81126 19009
rect 86040 18974 86092 18980
rect 81070 18935 81072 18944
rect 76116 18902 76144 18935
rect 81124 18935 81126 18944
rect 81072 18906 81124 18912
rect 76104 18896 76156 18902
rect 56046 18864 56102 18873
rect 56046 18799 56102 18808
rect 58162 18864 58218 18873
rect 58162 18799 58164 18808
rect 56060 18766 56088 18799
rect 58216 18799 58218 18808
rect 73710 18864 73766 18873
rect 76104 18838 76156 18844
rect 73710 18799 73712 18808
rect 58164 18770 58216 18776
rect 73764 18799 73766 18808
rect 73712 18770 73764 18776
rect 56048 18760 56100 18766
rect 56048 18702 56100 18708
rect 106094 18592 106150 18601
rect 106094 18527 106096 18536
rect 106148 18527 106150 18536
rect 108670 18592 108726 18601
rect 108670 18527 108726 18536
rect 106096 18498 106148 18504
rect 108684 18494 108712 18527
rect 108672 18488 108724 18494
rect 108672 18430 108724 18436
rect 113454 18456 113510 18465
rect 113454 18391 113456 18400
rect 113508 18391 113510 18400
rect 113456 18362 113508 18368
rect 62028 17944 62080 17950
rect 59542 17912 59598 17921
rect 59542 17847 59598 17856
rect 60462 17912 60518 17921
rect 60462 17847 60464 17856
rect 55956 17808 56008 17814
rect 55956 17750 56008 17756
rect 56508 17808 56560 17814
rect 56508 17750 56560 17756
rect 53840 17740 53892 17746
rect 53840 17682 53892 17688
rect 53852 17649 53880 17682
rect 53838 17640 53894 17649
rect 53472 17604 53524 17610
rect 53838 17575 53894 17584
rect 53472 17546 53524 17552
rect 56520 16862 56548 17750
rect 57886 17368 57942 17377
rect 57886 17303 57942 17312
rect 56508 16856 56560 16862
rect 56508 16798 56560 16804
rect 57900 16794 57928 17303
rect 59556 16930 59584 17847
rect 60516 17847 60518 17856
rect 62026 17912 62028 17921
rect 62080 17912 62082 17921
rect 62026 17847 62082 17856
rect 64694 17912 64750 17921
rect 64694 17847 64696 17856
rect 60464 17818 60516 17824
rect 64748 17847 64750 17856
rect 66166 17912 66222 17921
rect 66166 17847 66222 17856
rect 67638 17912 67694 17921
rect 67638 17847 67694 17856
rect 71778 17912 71834 17921
rect 71778 17847 71834 17856
rect 73158 17912 73214 17921
rect 73158 17847 73214 17856
rect 78586 17912 78642 17921
rect 78586 17847 78642 17856
rect 125966 17912 126022 17921
rect 125966 17847 126022 17856
rect 64696 17818 64748 17824
rect 60476 17474 60504 17818
rect 66180 17814 66208 17847
rect 66168 17808 66220 17814
rect 66168 17750 66220 17756
rect 67652 17542 67680 17847
rect 68928 17740 68980 17746
rect 68928 17682 68980 17688
rect 68940 17649 68968 17682
rect 68190 17640 68246 17649
rect 68190 17575 68246 17584
rect 68926 17640 68982 17649
rect 68926 17575 68982 17584
rect 70398 17640 70454 17649
rect 71792 17610 71820 17847
rect 70398 17575 70454 17584
rect 71780 17604 71832 17610
rect 67640 17536 67692 17542
rect 67640 17478 67692 17484
rect 60464 17468 60516 17474
rect 60464 17410 60516 17416
rect 67640 17400 67692 17406
rect 65062 17368 65118 17377
rect 65062 17303 65118 17312
rect 66258 17368 66314 17377
rect 66258 17303 66260 17312
rect 65076 17270 65104 17303
rect 66312 17303 66314 17312
rect 67638 17368 67640 17377
rect 68204 17377 68232 17575
rect 69662 17504 69718 17513
rect 69662 17439 69718 17448
rect 69676 17406 69704 17439
rect 69664 17400 69716 17406
rect 67692 17368 67694 17377
rect 67638 17303 67694 17312
rect 68190 17368 68246 17377
rect 69664 17342 69716 17348
rect 68190 17303 68246 17312
rect 66260 17274 66312 17280
rect 65064 17264 65116 17270
rect 60738 17232 60794 17241
rect 60738 17167 60794 17176
rect 62118 17232 62174 17241
rect 62118 17167 62174 17176
rect 63498 17232 63554 17241
rect 65064 17206 65116 17212
rect 69018 17232 69074 17241
rect 63498 17167 63500 17176
rect 60752 17066 60780 17167
rect 62132 17134 62160 17167
rect 63552 17167 63554 17176
rect 69018 17167 69074 17176
rect 63500 17138 63552 17144
rect 62120 17128 62172 17134
rect 62120 17070 62172 17076
rect 60740 17060 60792 17066
rect 60740 17002 60792 17008
rect 69032 16998 69060 17167
rect 69020 16992 69072 16998
rect 69020 16934 69072 16940
rect 59544 16924 59596 16930
rect 59544 16866 59596 16872
rect 57888 16788 57940 16794
rect 57888 16730 57940 16736
rect 70412 16726 70440 17575
rect 71780 17546 71832 17552
rect 71686 17232 71742 17241
rect 71686 17167 71688 17176
rect 71740 17167 71742 17176
rect 71688 17138 71740 17144
rect 73172 16862 73200 17847
rect 78600 17678 78628 17847
rect 78588 17672 78640 17678
rect 78588 17614 78640 17620
rect 83830 17640 83886 17649
rect 83830 17575 83886 17584
rect 83844 17542 83872 17575
rect 83832 17536 83884 17542
rect 75918 17504 75974 17513
rect 75918 17439 75974 17448
rect 78678 17504 78734 17513
rect 83832 17478 83884 17484
rect 88246 17504 88302 17513
rect 78678 17439 78680 17448
rect 75932 17406 75960 17439
rect 78732 17439 78734 17448
rect 88246 17439 88248 17448
rect 78680 17410 78732 17416
rect 88300 17439 88302 17448
rect 93582 17504 93638 17513
rect 93582 17439 93638 17448
rect 88248 17410 88300 17416
rect 93596 17406 93624 17439
rect 75920 17400 75972 17406
rect 75920 17342 75972 17348
rect 93584 17400 93636 17406
rect 93584 17342 93636 17348
rect 99286 17368 99342 17377
rect 99286 17303 99288 17312
rect 99340 17303 99342 17312
rect 111706 17368 111762 17377
rect 111706 17303 111762 17312
rect 99288 17274 99340 17280
rect 111720 17270 111748 17303
rect 111708 17264 111760 17270
rect 74814 17232 74870 17241
rect 111708 17206 111760 17212
rect 74814 17167 74870 17176
rect 73160 16856 73212 16862
rect 73160 16798 73212 16804
rect 74828 16794 74856 17167
rect 77298 16960 77354 16969
rect 77298 16895 77300 16904
rect 77352 16895 77354 16904
rect 77300 16866 77352 16872
rect 74816 16788 74868 16794
rect 74816 16730 74868 16736
rect 52368 16720 52420 16726
rect 52368 16662 52420 16668
rect 70400 16720 70452 16726
rect 70400 16662 70452 16668
rect 125980 16590 126008 17847
rect 157996 17270 158024 454990
rect 158076 450968 158128 450974
rect 158076 450910 158128 450916
rect 158088 107234 158116 450910
rect 158168 450016 158220 450022
rect 158168 449958 158220 449964
rect 158180 107370 158208 449958
rect 158732 189281 158760 579119
rect 159376 479602 159404 586910
rect 159468 489326 159496 587046
rect 159456 489320 159508 489326
rect 159456 489262 159508 489268
rect 159364 479596 159416 479602
rect 159364 479538 159416 479544
rect 162136 456210 162164 587318
rect 162216 586628 162268 586634
rect 162216 586570 162268 586576
rect 162228 472870 162256 586570
rect 162216 472864 162268 472870
rect 162216 472806 162268 472812
rect 163516 459066 163544 700606
rect 166264 700392 166316 700398
rect 166264 700334 166316 700340
rect 163596 586696 163648 586702
rect 163596 586638 163648 586644
rect 163608 483886 163636 586638
rect 163596 483880 163648 483886
rect 163596 483822 163648 483828
rect 166276 471442 166304 700334
rect 166356 586832 166408 586838
rect 166356 586774 166408 586780
rect 166264 471436 166316 471442
rect 166264 471378 166316 471384
rect 166368 471374 166396 586774
rect 167644 586560 167696 586566
rect 167644 586502 167696 586508
rect 166356 471368 166408 471374
rect 166356 471310 166408 471316
rect 167656 468586 167684 586502
rect 167644 468580 167696 468586
rect 167644 468522 167696 468528
rect 169772 461854 169800 702406
rect 175924 700596 175976 700602
rect 175924 700538 175976 700544
rect 174544 683188 174596 683194
rect 174544 683130 174596 683136
rect 174556 500546 174584 683130
rect 175936 500682 175964 700538
rect 191104 700528 191156 700534
rect 191104 700470 191156 700476
rect 180064 700460 180116 700466
rect 180064 700402 180116 700408
rect 175924 500676 175976 500682
rect 175924 500618 175976 500624
rect 174544 500540 174596 500546
rect 174544 500482 174596 500488
rect 173346 463040 173402 463049
rect 173346 462975 173402 462984
rect 173162 462768 173218 462777
rect 173162 462703 173218 462712
rect 170402 462632 170458 462641
rect 170402 462567 170458 462576
rect 169760 461848 169812 461854
rect 169760 461790 169812 461796
rect 163504 459060 163556 459066
rect 163504 459002 163556 459008
rect 162124 456204 162176 456210
rect 162124 456146 162176 456152
rect 165620 246356 165672 246362
rect 165620 246298 165672 246304
rect 161480 244928 161532 244934
rect 161480 244870 161532 244876
rect 158718 189272 158774 189281
rect 158718 189207 158774 189216
rect 158168 107364 158220 107370
rect 158168 107306 158220 107312
rect 158076 107228 158128 107234
rect 158076 107170 158128 107176
rect 158732 99249 158760 189207
rect 158718 99240 158774 99249
rect 158718 99175 158774 99184
rect 158902 99240 158958 99249
rect 158902 99175 158958 99184
rect 158916 98666 158944 99175
rect 158904 98660 158956 98666
rect 158904 98602 158956 98608
rect 157984 17264 158036 17270
rect 157984 17206 158036 17212
rect 125968 16584 126020 16590
rect 161492 16574 161520 244870
rect 165632 16574 165660 246298
rect 170416 17202 170444 462567
rect 172520 243568 172572 243574
rect 172520 243510 172572 243516
rect 170496 98660 170548 98666
rect 170496 98602 170548 98608
rect 170508 57934 170536 98602
rect 170496 57928 170548 57934
rect 170496 57870 170548 57876
rect 170404 17196 170456 17202
rect 170404 17138 170456 17144
rect 172532 16574 172560 243510
rect 173176 17814 173204 462703
rect 173254 461272 173310 461281
rect 173254 461207 173310 461216
rect 173164 17808 173216 17814
rect 173164 17750 173216 17756
rect 173268 17746 173296 461207
rect 173360 17950 173388 462975
rect 175922 462496 175978 462505
rect 175922 462431 175978 462440
rect 173530 462360 173586 462369
rect 173530 462295 173586 462304
rect 173440 461032 173492 461038
rect 173440 460974 173492 460980
rect 173348 17944 173400 17950
rect 173348 17886 173400 17892
rect 173452 17882 173480 460974
rect 173544 19145 173572 462295
rect 173624 461100 173676 461106
rect 173624 461042 173676 461048
rect 173530 19136 173586 19145
rect 173530 19071 173586 19080
rect 173636 18766 173664 461042
rect 173714 461000 173770 461009
rect 173714 460935 173770 460944
rect 173728 19281 173756 460935
rect 173806 456240 173862 456249
rect 173806 456175 173862 456184
rect 173714 19272 173770 19281
rect 173714 19207 173770 19216
rect 173624 18760 173676 18766
rect 173624 18702 173676 18708
rect 173820 18698 173848 456175
rect 174544 247920 174596 247926
rect 174544 247862 174596 247868
rect 173808 18692 173860 18698
rect 173808 18634 173860 18640
rect 173440 17876 173492 17882
rect 173440 17818 173492 17824
rect 173256 17740 173308 17746
rect 173256 17682 173308 17688
rect 161492 16546 162072 16574
rect 165632 16546 166120 16574
rect 172532 16546 172744 16574
rect 125968 16526 126020 16532
rect 130568 15904 130620 15910
rect 130568 15846 130620 15852
rect 126980 14476 127032 14482
rect 126980 14418 127032 14424
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 125876 4820 125928 4826
rect 125876 4762 125928 4768
rect 125888 480 125916 4762
rect 126992 480 127020 14418
rect 128176 10328 128228 10334
rect 128176 10270 128228 10276
rect 128188 480 128216 10270
rect 130580 480 130608 15846
rect 158904 7608 158956 7614
rect 158904 7550 158956 7556
rect 155408 3868 155460 3874
rect 155408 3810 155460 3816
rect 151820 3800 151872 3806
rect 151820 3742 151872 3748
rect 144736 3732 144788 3738
rect 144736 3674 144788 3680
rect 137652 3664 137704 3670
rect 137652 3606 137704 3612
rect 134156 3596 134208 3602
rect 134156 3538 134208 3544
rect 134168 480 134196 3538
rect 137664 480 137692 3606
rect 141240 3460 141292 3466
rect 141240 3402 141292 3408
rect 141252 480 141280 3402
rect 144748 480 144776 3674
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148336 480 148364 3470
rect 151832 480 151860 3742
rect 155420 480 155448 3810
rect 158916 480 158944 7550
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 166092 480 166120 16546
rect 169576 6180 169628 6186
rect 169576 6122 169628 6128
rect 169588 480 169616 6122
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 174556 3806 174584 247862
rect 175832 247852 175884 247858
rect 175832 247794 175884 247800
rect 175844 3874 175872 247794
rect 175936 18494 175964 462431
rect 176106 461136 176162 461145
rect 176106 461071 176162 461080
rect 176014 459776 176070 459785
rect 176014 459711 176070 459720
rect 175924 18488 175976 18494
rect 175924 18430 175976 18436
rect 176028 17338 176056 459711
rect 176120 18426 176148 461071
rect 179326 460320 179382 460329
rect 179326 460255 179382 460264
rect 179142 460048 179198 460057
rect 179142 459983 179198 459992
rect 178590 459912 178646 459921
rect 178590 459847 178646 459856
rect 176198 459640 176254 459649
rect 176198 459575 176254 459584
rect 176212 19310 176240 459575
rect 176290 458688 176346 458697
rect 176290 458623 176346 458632
rect 176200 19304 176252 19310
rect 176200 19246 176252 19252
rect 176304 19242 176332 458623
rect 176474 458552 176530 458561
rect 176474 458487 176530 458496
rect 176382 457600 176438 457609
rect 176382 457535 176438 457544
rect 176292 19236 176344 19242
rect 176292 19178 176344 19184
rect 176396 18630 176424 457535
rect 176384 18624 176436 18630
rect 176384 18566 176436 18572
rect 176488 18562 176516 458487
rect 176566 452976 176622 452985
rect 176566 452911 176622 452920
rect 176580 19174 176608 452911
rect 177304 451852 177356 451858
rect 177304 451794 177356 451800
rect 177316 346390 177344 451794
rect 177304 346384 177356 346390
rect 177304 346326 177356 346332
rect 176660 242208 176712 242214
rect 176660 242150 176712 242156
rect 176568 19168 176620 19174
rect 176568 19110 176620 19116
rect 176476 18556 176528 18562
rect 176476 18498 176528 18504
rect 176108 18420 176160 18426
rect 176108 18362 176160 18368
rect 176016 17332 176068 17338
rect 176016 17274 176068 17280
rect 175832 3868 175884 3874
rect 175832 3810 175884 3816
rect 174544 3800 174596 3806
rect 174544 3742 174596 3748
rect 176672 480 176700 242150
rect 178604 19106 178632 459847
rect 179052 459672 179104 459678
rect 179052 459614 179104 459620
rect 178776 459196 178828 459202
rect 178776 459138 178828 459144
rect 178684 458448 178736 458454
rect 178684 458390 178736 458396
rect 178592 19100 178644 19106
rect 178592 19042 178644 19048
rect 178696 17542 178724 458390
rect 178788 17678 178816 459138
rect 178958 458824 179014 458833
rect 178958 458759 179014 458768
rect 178868 458380 178920 458386
rect 178868 458322 178920 458328
rect 178776 17672 178828 17678
rect 178776 17614 178828 17620
rect 178684 17536 178736 17542
rect 178684 17478 178736 17484
rect 178880 17474 178908 458322
rect 178868 17468 178920 17474
rect 178868 17410 178920 17416
rect 178972 17406 179000 458759
rect 179064 18902 179092 459614
rect 179156 19038 179184 459983
rect 179236 247988 179288 247994
rect 179236 247930 179288 247936
rect 179144 19032 179196 19038
rect 179144 18974 179196 18980
rect 179052 18896 179104 18902
rect 179052 18838 179104 18844
rect 178960 17400 179012 17406
rect 178960 17342 179012 17348
rect 179248 3738 179276 247930
rect 179340 18970 179368 460255
rect 180076 459134 180104 700402
rect 187608 464500 187660 464506
rect 187608 464442 187660 464448
rect 186872 464432 186924 464438
rect 186872 464374 186924 464380
rect 186780 464092 186832 464098
rect 186780 464034 186832 464040
rect 183468 464024 183520 464030
rect 183468 463966 183520 463972
rect 181444 459808 181496 459814
rect 181444 459750 181496 459756
rect 180064 459128 180116 459134
rect 180064 459070 180116 459076
rect 181352 454980 181404 454986
rect 181352 454922 181404 454928
rect 181364 293962 181392 454922
rect 181352 293956 181404 293962
rect 181352 293898 181404 293904
rect 181352 248056 181404 248062
rect 181352 247998 181404 248004
rect 179420 239420 179472 239426
rect 179420 239362 179472 239368
rect 179328 18964 179380 18970
rect 179328 18906 179380 18912
rect 179432 16574 179460 239362
rect 179432 16546 180288 16574
rect 179236 3732 179288 3738
rect 179236 3674 179288 3680
rect 180260 480 180288 16546
rect 181364 3602 181392 247998
rect 181456 17785 181484 459750
rect 181720 459740 181772 459746
rect 181720 459682 181772 459688
rect 181628 459604 181680 459610
rect 181628 459546 181680 459552
rect 181536 459264 181588 459270
rect 181536 459206 181588 459212
rect 181548 18834 181576 459206
rect 181640 107098 181668 459546
rect 181732 108594 181760 459682
rect 181904 458516 181956 458522
rect 181904 458458 181956 458464
rect 181810 457056 181866 457065
rect 181810 456991 181866 457000
rect 181720 108588 181772 108594
rect 181720 108530 181772 108536
rect 181824 107166 181852 456991
rect 181916 108662 181944 458458
rect 181996 456408 182048 456414
rect 181996 456350 182048 456356
rect 181904 108656 181956 108662
rect 181904 108598 181956 108604
rect 182008 108526 182036 456350
rect 183376 456340 183428 456346
rect 183376 456282 183428 456288
rect 182824 450628 182876 450634
rect 182824 450570 182876 450576
rect 182088 450220 182140 450226
rect 182088 450162 182140 450168
rect 181996 108520 182048 108526
rect 181996 108462 182048 108468
rect 181812 107160 181864 107166
rect 181812 107102 181864 107108
rect 181628 107092 181680 107098
rect 181628 107034 181680 107040
rect 182100 106729 182128 450162
rect 182836 202842 182864 450570
rect 182916 248124 182968 248130
rect 182916 248066 182968 248072
rect 182824 202836 182876 202842
rect 182824 202778 182876 202784
rect 182086 106720 182142 106729
rect 182086 106655 182142 106664
rect 181536 18828 181588 18834
rect 181536 18770 181588 18776
rect 181442 17776 181498 17785
rect 181442 17711 181498 17720
rect 182928 3670 182956 248066
rect 183388 17678 183416 456282
rect 183480 17746 183508 463966
rect 186228 463956 186280 463962
rect 186228 463898 186280 463904
rect 184848 463888 184900 463894
rect 184848 463830 184900 463836
rect 184756 458720 184808 458726
rect 184756 458662 184808 458668
rect 184204 457088 184256 457094
rect 184204 457030 184256 457036
rect 184020 454912 184072 454918
rect 184020 454854 184072 454860
rect 184032 358766 184060 454854
rect 184112 450356 184164 450362
rect 184112 450298 184164 450304
rect 184020 358760 184072 358766
rect 184020 358702 184072 358708
rect 184124 108458 184152 450298
rect 184216 108798 184244 457030
rect 184296 457020 184348 457026
rect 184296 456962 184348 456968
rect 184308 108934 184336 456962
rect 184480 455864 184532 455870
rect 184480 455806 184532 455812
rect 184388 455796 184440 455802
rect 184388 455738 184440 455744
rect 184400 109002 184428 455738
rect 184388 108996 184440 109002
rect 184388 108938 184440 108944
rect 184296 108928 184348 108934
rect 184296 108870 184348 108876
rect 184492 108866 184520 455806
rect 184570 451616 184626 451625
rect 184570 451551 184626 451560
rect 184480 108860 184532 108866
rect 184480 108802 184532 108808
rect 184204 108792 184256 108798
rect 184204 108734 184256 108740
rect 184112 108452 184164 108458
rect 184112 108394 184164 108400
rect 184584 108390 184612 451551
rect 184662 450120 184718 450129
rect 184662 450055 184718 450064
rect 184676 108730 184704 450055
rect 184664 108724 184716 108730
rect 184664 108666 184716 108672
rect 184572 108384 184624 108390
rect 184572 108326 184624 108332
rect 183560 102808 183612 102814
rect 183560 102750 183612 102756
rect 183468 17740 183520 17746
rect 183468 17682 183520 17688
rect 183376 17672 183428 17678
rect 183376 17614 183428 17620
rect 183572 16574 183600 102750
rect 184768 17474 184796 458662
rect 184756 17468 184808 17474
rect 184756 17410 184808 17416
rect 184860 17270 184888 463830
rect 186136 463820 186188 463826
rect 186136 463762 186188 463768
rect 185860 461372 185912 461378
rect 185860 461314 185912 461320
rect 185768 461168 185820 461174
rect 185768 461110 185820 461116
rect 185400 453076 185452 453082
rect 185400 453018 185452 453024
rect 185412 241466 185440 453018
rect 185492 452804 185544 452810
rect 185492 452746 185544 452752
rect 185400 241460 185452 241466
rect 185400 241402 185452 241408
rect 185504 18873 185532 452746
rect 185584 452736 185636 452742
rect 185584 452678 185636 452684
rect 185596 19145 185624 452678
rect 185676 451784 185728 451790
rect 185676 451726 185728 451732
rect 185582 19136 185638 19145
rect 185582 19071 185638 19080
rect 185490 18864 185546 18873
rect 185490 18799 185546 18808
rect 185688 17950 185716 451726
rect 185780 18630 185808 461110
rect 185872 18698 185900 461314
rect 185952 459944 186004 459950
rect 185952 459886 186004 459892
rect 185860 18692 185912 18698
rect 185860 18634 185912 18640
rect 185768 18624 185820 18630
rect 185768 18566 185820 18572
rect 185676 17944 185728 17950
rect 185676 17886 185728 17892
rect 185964 17542 185992 459886
rect 186044 459876 186096 459882
rect 186044 459818 186096 459824
rect 185952 17536 186004 17542
rect 185952 17478 186004 17484
rect 186056 17406 186084 459818
rect 186044 17400 186096 17406
rect 186044 17342 186096 17348
rect 186148 17338 186176 463762
rect 186136 17332 186188 17338
rect 186136 17274 186188 17280
rect 184848 17264 184900 17270
rect 184848 17206 184900 17212
rect 186240 17202 186268 463898
rect 186792 394777 186820 464034
rect 186778 394768 186834 394777
rect 186778 394703 186834 394712
rect 186884 250510 186912 464374
rect 186964 457224 187016 457230
rect 186964 457166 187016 457172
rect 186872 250504 186924 250510
rect 186872 250446 186924 250452
rect 186318 247616 186374 247625
rect 186318 247551 186374 247560
rect 186228 17196 186280 17202
rect 186228 17138 186280 17144
rect 186332 16574 186360 247551
rect 186976 107574 187004 457166
rect 187056 457156 187108 457162
rect 187056 457098 187108 457104
rect 186964 107568 187016 107574
rect 186964 107510 187016 107516
rect 187068 107438 187096 457098
rect 187240 456272 187292 456278
rect 187240 456214 187292 456220
rect 187148 456000 187200 456006
rect 187148 455942 187200 455948
rect 187160 107506 187188 455942
rect 187252 108322 187280 456214
rect 187516 454640 187568 454646
rect 187516 454582 187568 454588
rect 187330 453384 187386 453393
rect 187330 453319 187386 453328
rect 187344 215286 187372 453319
rect 187424 450424 187476 450430
rect 187424 450366 187476 450372
rect 187332 215280 187384 215286
rect 187332 215222 187384 215228
rect 187240 108316 187292 108322
rect 187240 108258 187292 108264
rect 187148 107500 187200 107506
rect 187148 107442 187200 107448
rect 187056 107432 187108 107438
rect 187056 107374 187108 107380
rect 187436 17377 187464 450366
rect 187528 18970 187556 454582
rect 187516 18964 187568 18970
rect 187516 18906 187568 18912
rect 187620 17882 187648 464442
rect 188988 464296 189040 464302
rect 188988 464238 189040 464244
rect 188160 464160 188212 464166
rect 188160 464102 188212 464108
rect 188068 452940 188120 452946
rect 188068 452882 188120 452888
rect 188080 446486 188108 452882
rect 188068 446480 188120 446486
rect 188068 446422 188120 446428
rect 188172 369073 188200 464102
rect 188620 458992 188672 458998
rect 188620 458934 188672 458940
rect 188436 453008 188488 453014
rect 188436 452950 188488 452956
rect 188342 451752 188398 451761
rect 188342 451687 188398 451696
rect 188252 450696 188304 450702
rect 188252 450638 188304 450644
rect 188158 369064 188214 369073
rect 188158 368999 188214 369008
rect 188264 320142 188292 450638
rect 188252 320136 188304 320142
rect 188252 320078 188304 320084
rect 188356 19009 188384 451687
rect 188448 447982 188476 452950
rect 188528 452872 188580 452878
rect 188528 452814 188580 452820
rect 188436 447976 188488 447982
rect 188436 447918 188488 447924
rect 188436 446480 188488 446486
rect 188436 446422 188488 446428
rect 188342 19000 188398 19009
rect 188342 18935 188398 18944
rect 188448 18494 188476 446422
rect 188540 19174 188568 452814
rect 188632 451314 188660 458934
rect 188712 454844 188764 454850
rect 188712 454786 188764 454792
rect 188620 451308 188672 451314
rect 188620 451250 188672 451256
rect 188620 447976 188672 447982
rect 188620 447918 188672 447924
rect 188528 19168 188580 19174
rect 188528 19110 188580 19116
rect 188632 19106 188660 447918
rect 188620 19100 188672 19106
rect 188620 19042 188672 19048
rect 188724 18562 188752 454786
rect 188804 454776 188856 454782
rect 188804 454718 188856 454724
rect 188816 19310 188844 454718
rect 188896 451580 188948 451586
rect 188896 451522 188948 451528
rect 188908 451489 188936 451522
rect 188894 451480 188950 451489
rect 188894 451415 188950 451424
rect 188896 451308 188948 451314
rect 188896 451250 188948 451256
rect 188804 19304 188856 19310
rect 188804 19246 188856 19252
rect 188908 18737 188936 451250
rect 189000 19378 189028 464238
rect 191116 461922 191144 700470
rect 192484 700324 192536 700330
rect 192484 700266 192536 700272
rect 191472 464228 191524 464234
rect 191472 464170 191524 464176
rect 191104 461916 191156 461922
rect 191104 461858 191156 461864
rect 189540 461304 189592 461310
rect 189540 461246 189592 461252
rect 189552 397458 189580 461246
rect 190368 461236 190420 461242
rect 190368 461178 190420 461184
rect 190276 458788 190328 458794
rect 190276 458730 190328 458736
rect 190090 452024 190146 452033
rect 189632 451988 189684 451994
rect 190090 451959 190146 451968
rect 189632 451930 189684 451936
rect 189540 397452 189592 397458
rect 189540 397394 189592 397400
rect 189644 267714 189672 451930
rect 189998 451888 190054 451897
rect 189998 451823 190054 451832
rect 189816 450492 189868 450498
rect 189816 450434 189868 450440
rect 189724 449540 189776 449546
rect 189724 449482 189776 449488
rect 189632 267708 189684 267714
rect 189632 267650 189684 267656
rect 189736 53718 189764 449482
rect 189828 53786 189856 450434
rect 189908 449608 189960 449614
rect 189908 449550 189960 449556
rect 189816 53780 189868 53786
rect 189816 53722 189868 53728
rect 189724 53712 189776 53718
rect 189724 53654 189776 53660
rect 189920 52426 189948 449550
rect 189908 52420 189960 52426
rect 189908 52362 189960 52368
rect 190012 51066 190040 451823
rect 190000 51060 190052 51066
rect 190000 51002 190052 51008
rect 190104 48278 190132 451959
rect 190184 449676 190236 449682
rect 190184 449618 190236 449624
rect 190092 48272 190144 48278
rect 190092 48214 190144 48220
rect 188988 19372 189040 19378
rect 188988 19314 189040 19320
rect 190196 18902 190224 449618
rect 190288 19242 190316 458730
rect 190276 19236 190328 19242
rect 190276 19178 190328 19184
rect 190184 18896 190236 18902
rect 190184 18838 190236 18844
rect 190380 18834 190408 461178
rect 191012 453144 191064 453150
rect 191012 453086 191064 453092
rect 190920 452056 190972 452062
rect 190920 451998 190972 452004
rect 190826 398848 190882 398857
rect 190826 398783 190828 398792
rect 190880 398783 190882 398792
rect 190828 398754 190880 398760
rect 190828 397452 190880 397458
rect 190828 397394 190880 397400
rect 190840 397361 190868 397394
rect 190826 397352 190882 397361
rect 190826 397287 190882 397296
rect 190826 372600 190882 372609
rect 190826 372535 190828 372544
rect 190880 372535 190882 372544
rect 190828 372506 190880 372512
rect 190932 306338 190960 451998
rect 190920 306332 190972 306338
rect 190920 306274 190972 306280
rect 191024 258074 191052 453086
rect 191380 452124 191432 452130
rect 191380 452066 191432 452072
rect 191288 451920 191340 451926
rect 191288 451862 191340 451868
rect 191104 450764 191156 450770
rect 191104 450706 191156 450712
rect 191116 398857 191144 450706
rect 191196 450288 191248 450294
rect 191196 450230 191248 450236
rect 191102 398848 191158 398857
rect 191102 398783 191158 398792
rect 191102 397352 191158 397361
rect 191102 397287 191158 397296
rect 190932 258046 191052 258074
rect 190932 255270 190960 258046
rect 190920 255264 190972 255270
rect 190920 255206 190972 255212
rect 190368 18828 190420 18834
rect 190368 18770 190420 18776
rect 188894 18728 188950 18737
rect 188894 18663 188950 18672
rect 188712 18556 188764 18562
rect 188712 18498 188764 18504
rect 188436 18488 188488 18494
rect 188436 18430 188488 18436
rect 187608 17876 187660 17882
rect 187608 17818 187660 17824
rect 187422 17368 187478 17377
rect 187422 17303 187478 17312
rect 191116 17066 191144 397287
rect 191208 107642 191236 450230
rect 191300 217326 191328 451862
rect 191392 372609 191420 452066
rect 191484 419665 191512 464170
rect 192496 461990 192524 700266
rect 199936 682644 199988 682650
rect 199936 682586 199988 682592
rect 196624 682576 196676 682582
rect 196624 682518 196676 682524
rect 196532 682508 196584 682514
rect 196532 682450 196584 682456
rect 195060 682440 195112 682446
rect 195060 682382 195112 682388
rect 194416 680672 194468 680678
rect 194416 680614 194468 680620
rect 193036 680604 193088 680610
rect 193036 680546 193088 680552
rect 193048 499050 193076 680546
rect 193128 680536 193180 680542
rect 193128 680478 193180 680484
rect 193036 499044 193088 499050
rect 193036 498986 193088 498992
rect 193140 494970 193168 680478
rect 194428 499118 194456 680614
rect 194508 680468 194560 680474
rect 194508 680410 194560 680416
rect 194416 499112 194468 499118
rect 194416 499054 194468 499060
rect 194520 495038 194548 680410
rect 195072 500410 195100 682382
rect 195888 682032 195940 682038
rect 195888 681974 195940 681980
rect 195520 680944 195572 680950
rect 195520 680886 195572 680892
rect 195428 680400 195480 680406
rect 195428 680342 195480 680348
rect 195152 679652 195204 679658
rect 195152 679594 195204 679600
rect 195060 500404 195112 500410
rect 195060 500346 195112 500352
rect 195164 497826 195192 679594
rect 195242 679416 195298 679425
rect 195242 679351 195298 679360
rect 195256 498030 195284 679351
rect 195334 679280 195390 679289
rect 195334 679215 195390 679224
rect 195244 498024 195296 498030
rect 195244 497966 195296 497972
rect 195152 497820 195204 497826
rect 195152 497762 195204 497768
rect 195348 497554 195376 679215
rect 195440 498137 195468 680342
rect 195426 498128 195482 498137
rect 195532 498098 195560 680886
rect 195704 679584 195756 679590
rect 195704 679526 195756 679532
rect 195612 679516 195664 679522
rect 195612 679458 195664 679464
rect 195426 498063 195482 498072
rect 195520 498092 195572 498098
rect 195520 498034 195572 498040
rect 195336 497548 195388 497554
rect 195336 497490 195388 497496
rect 194508 495032 194560 495038
rect 194508 494974 194560 494980
rect 193128 494964 193180 494970
rect 193128 494906 193180 494912
rect 195624 466138 195652 679458
rect 195716 466274 195744 679526
rect 195796 679448 195848 679454
rect 195796 679390 195848 679396
rect 195704 466268 195756 466274
rect 195704 466210 195756 466216
rect 195612 466132 195664 466138
rect 195612 466074 195664 466080
rect 195808 465934 195836 679390
rect 195796 465928 195848 465934
rect 195796 465870 195848 465876
rect 195900 463418 195928 681974
rect 196438 678328 196494 678337
rect 196438 678263 196494 678272
rect 196452 498166 196480 678263
rect 196544 500614 196572 682450
rect 196532 500608 196584 500614
rect 196532 500550 196584 500556
rect 196636 500274 196664 682518
rect 196716 682372 196768 682378
rect 196716 682314 196768 682320
rect 196728 500478 196756 682314
rect 199660 682304 199712 682310
rect 199660 682246 199712 682252
rect 196806 682136 196862 682145
rect 196806 682071 196862 682080
rect 199384 682100 199436 682106
rect 196716 500472 196768 500478
rect 196716 500414 196768 500420
rect 196820 500342 196848 682071
rect 199384 682042 199436 682048
rect 198648 681828 198700 681834
rect 198648 681770 198700 681776
rect 197084 680876 197136 680882
rect 197084 680818 197136 680824
rect 196990 679688 197046 679697
rect 196990 679623 197046 679632
rect 196898 679144 196954 679153
rect 196898 679079 196954 679088
rect 196808 500336 196860 500342
rect 196808 500278 196860 500284
rect 196624 500268 196676 500274
rect 196624 500210 196676 500216
rect 196440 498160 196492 498166
rect 196440 498102 196492 498108
rect 196912 497622 196940 679079
rect 197004 497690 197032 679623
rect 197096 497894 197124 680818
rect 197176 680808 197228 680814
rect 197176 680750 197228 680756
rect 197084 497888 197136 497894
rect 197084 497830 197136 497836
rect 196992 497684 197044 497690
rect 196992 497626 197044 497632
rect 196900 497616 196952 497622
rect 196900 497558 196952 497564
rect 197188 497418 197216 680750
rect 198464 680740 198516 680746
rect 198464 680682 198516 680688
rect 197268 679448 197320 679454
rect 197268 679390 197320 679396
rect 197176 497412 197228 497418
rect 197176 497354 197228 497360
rect 197280 468654 197308 679390
rect 197820 584996 197872 585002
rect 197820 584938 197872 584944
rect 197268 468648 197320 468654
rect 197268 468590 197320 468596
rect 197832 466041 197860 584938
rect 197912 584928 197964 584934
rect 197912 584870 197964 584876
rect 197818 466032 197874 466041
rect 197818 465967 197874 465976
rect 197924 465866 197952 584870
rect 198188 584860 198240 584866
rect 198188 584802 198240 584808
rect 198004 584656 198056 584662
rect 198004 584598 198056 584604
rect 197912 465860 197964 465866
rect 197912 465802 197964 465808
rect 195888 463412 195940 463418
rect 195888 463354 195940 463360
rect 192484 461984 192536 461990
rect 192484 461926 192536 461932
rect 191748 461440 191800 461446
rect 191748 461382 191800 461388
rect 191656 457292 191708 457298
rect 191656 457234 191708 457240
rect 191564 452668 191616 452674
rect 191564 452610 191616 452616
rect 191470 419656 191526 419665
rect 191470 419591 191526 419600
rect 191470 397352 191526 397361
rect 191470 397287 191526 397296
rect 191378 372600 191434 372609
rect 191378 372535 191434 372544
rect 191378 369880 191434 369889
rect 191378 369815 191434 369824
rect 191288 217320 191340 217326
rect 191288 217262 191340 217268
rect 191196 107636 191248 107642
rect 191196 107578 191248 107584
rect 191392 17513 191420 369815
rect 191484 17814 191512 397287
rect 191576 56574 191604 452610
rect 191564 56568 191616 56574
rect 191564 56510 191616 56516
rect 191668 18766 191696 457234
rect 191760 19038 191788 461382
rect 198016 460562 198044 584598
rect 198096 584588 198148 584594
rect 198096 584530 198148 584536
rect 198108 460630 198136 584530
rect 198096 460624 198148 460630
rect 198096 460566 198148 460572
rect 198004 460556 198056 460562
rect 198004 460498 198056 460504
rect 198200 460358 198228 584802
rect 198280 584792 198332 584798
rect 198280 584734 198332 584740
rect 198292 460426 198320 584734
rect 198372 584724 198424 584730
rect 198372 584666 198424 584672
rect 198384 460494 198412 584666
rect 198476 497729 198504 680682
rect 198556 679312 198608 679318
rect 198556 679254 198608 679260
rect 198462 497720 198518 497729
rect 198462 497655 198518 497664
rect 198568 466002 198596 679254
rect 198660 466410 198688 681770
rect 199290 679824 199346 679833
rect 199290 679759 199346 679768
rect 199198 678192 199254 678201
rect 199198 678127 199254 678136
rect 199212 497962 199240 678127
rect 199200 497956 199252 497962
rect 199200 497898 199252 497904
rect 198648 466404 198700 466410
rect 198648 466346 198700 466352
rect 198556 465996 198608 466002
rect 198556 465938 198608 465944
rect 199304 465594 199332 679759
rect 199396 466206 199424 682042
rect 199568 681964 199620 681970
rect 199568 681906 199620 681912
rect 199474 679552 199530 679561
rect 199474 679487 199530 679496
rect 199384 466200 199436 466206
rect 199384 466142 199436 466148
rect 199292 465588 199344 465594
rect 199292 465530 199344 465536
rect 199488 462874 199516 679487
rect 199580 462942 199608 681906
rect 199672 463554 199700 682246
rect 199844 682236 199896 682242
rect 199844 682178 199896 682184
rect 199752 681896 199804 681902
rect 199752 681838 199804 681844
rect 199764 463690 199792 681838
rect 199752 463684 199804 463690
rect 199752 463626 199804 463632
rect 199660 463548 199712 463554
rect 199660 463490 199712 463496
rect 199856 463486 199884 682178
rect 199948 463622 199976 682586
rect 201222 682272 201278 682281
rect 201222 682207 201278 682216
rect 201130 682000 201186 682009
rect 201130 681935 201186 681944
rect 200028 681760 200080 681766
rect 200028 681702 200080 681708
rect 199936 463616 199988 463622
rect 199936 463558 199988 463564
rect 199844 463480 199896 463486
rect 199844 463422 199896 463428
rect 199568 462936 199620 462942
rect 199568 462878 199620 462884
rect 199476 462868 199528 462874
rect 199476 462810 199528 462816
rect 198740 460964 198792 460970
rect 198792 460912 199700 460934
rect 198740 460906 199700 460912
rect 198372 460488 198424 460494
rect 198372 460430 198424 460436
rect 198280 460420 198332 460426
rect 198280 460362 198332 460368
rect 198188 460352 198240 460358
rect 198188 460294 198240 460300
rect 197542 458416 197598 458425
rect 197542 458351 197598 458360
rect 195978 458280 196034 458289
rect 195978 458215 196034 458224
rect 195992 456794 196020 458215
rect 195992 456766 196388 456794
rect 196254 455560 196310 455569
rect 196254 455495 196310 455504
rect 194598 454200 194654 454209
rect 194598 454135 194654 454144
rect 193864 453212 193916 453218
rect 193864 453154 193916 453160
rect 193678 452704 193734 452713
rect 193678 452639 193734 452648
rect 193692 449956 193720 452639
rect 191840 449948 191892 449954
rect 191840 449890 191892 449896
rect 191852 422385 191880 449890
rect 193876 449886 193904 453154
rect 194506 450800 194562 450809
rect 194506 450735 194562 450744
rect 194520 450537 194548 450735
rect 194322 450528 194378 450537
rect 194322 450463 194378 450472
rect 194506 450528 194562 450537
rect 194506 450463 194562 450472
rect 194336 450265 194364 450463
rect 194138 450256 194194 450265
rect 194138 450191 194194 450200
rect 194322 450256 194378 450265
rect 194322 450191 194378 450200
rect 194152 449970 194180 450191
rect 194612 449970 194640 454135
rect 195520 451580 195572 451586
rect 195520 451522 195572 451528
rect 195150 451480 195206 451489
rect 195150 451415 195206 451424
rect 194152 449942 194442 449970
rect 194612 449942 194810 449970
rect 195164 449956 195192 451415
rect 195532 449956 195560 451522
rect 195886 451344 195942 451353
rect 195886 451279 195942 451288
rect 195900 449956 195928 451279
rect 196268 449956 196296 455495
rect 196360 449970 196388 456766
rect 197358 455696 197414 455705
rect 197358 455631 197414 455640
rect 196990 454064 197046 454073
rect 196990 453999 197046 454008
rect 196360 449942 196650 449970
rect 197004 449956 197032 453999
rect 197372 449956 197400 455631
rect 197556 449970 197584 458351
rect 198832 458312 198884 458318
rect 198832 458254 198884 458260
rect 198464 455456 198516 455462
rect 198464 455398 198516 455404
rect 198096 454096 198148 454102
rect 198096 454038 198148 454044
rect 197556 449942 197754 449970
rect 198108 449956 198136 454038
rect 198476 449956 198504 455398
rect 198844 449956 198872 458254
rect 199292 458244 199344 458250
rect 199292 458186 199344 458192
rect 199200 454436 199252 454442
rect 199200 454378 199252 454384
rect 199212 449956 199240 454378
rect 199304 449970 199332 458186
rect 199672 449970 199700 460906
rect 200040 460698 200068 681702
rect 200868 585138 201080 585154
rect 200856 585132 201080 585138
rect 200908 585126 201080 585132
rect 200856 585074 200908 585080
rect 200948 585064 201000 585070
rect 200948 585006 201000 585012
rect 200672 584520 200724 584526
rect 200672 584462 200724 584468
rect 200580 584452 200632 584458
rect 200580 584394 200632 584400
rect 200592 463350 200620 584394
rect 200580 463344 200632 463350
rect 200580 463286 200632 463292
rect 200684 463282 200712 584462
rect 200764 584384 200816 584390
rect 200764 584326 200816 584332
rect 200672 463276 200724 463282
rect 200672 463218 200724 463224
rect 200776 460934 200804 584326
rect 200856 584316 200908 584322
rect 200856 584258 200908 584264
rect 200868 461786 200896 584258
rect 200960 463214 200988 585006
rect 200948 463208 201000 463214
rect 200948 463150 201000 463156
rect 201052 463146 201080 585126
rect 201144 501673 201172 681935
rect 201130 501664 201186 501673
rect 201130 501599 201186 501608
rect 201236 497758 201264 682207
rect 201316 679176 201368 679182
rect 201316 679118 201368 679124
rect 201224 497752 201276 497758
rect 201224 497694 201276 497700
rect 201328 468722 201356 679118
rect 201408 679040 201460 679046
rect 201408 678982 201460 678988
rect 201316 468716 201368 468722
rect 201316 468658 201368 468664
rect 201420 465662 201448 678982
rect 201512 481098 201540 702986
rect 218992 700913 219020 703520
rect 218978 700904 219034 700913
rect 218978 700839 219034 700848
rect 235184 700466 235212 703520
rect 202144 700460 202196 700466
rect 202144 700402 202196 700408
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 202052 700324 202104 700330
rect 202052 700266 202104 700272
rect 201866 682816 201922 682825
rect 201866 682751 201922 682760
rect 201684 679856 201736 679862
rect 201684 679798 201736 679804
rect 201592 679244 201644 679250
rect 201592 679186 201644 679192
rect 201604 496262 201632 679186
rect 201696 679046 201724 679798
rect 201776 679312 201828 679318
rect 201776 679254 201828 679260
rect 201684 679040 201736 679046
rect 201684 678982 201736 678988
rect 201788 678910 201816 679254
rect 201776 678904 201828 678910
rect 201776 678846 201828 678852
rect 201880 669314 201908 682751
rect 201960 682168 202012 682174
rect 201960 682110 202012 682116
rect 201972 678366 202000 682110
rect 201960 678360 202012 678366
rect 201960 678302 202012 678308
rect 201880 669286 202000 669314
rect 201972 500750 202000 669286
rect 202064 501362 202092 700266
rect 202052 501356 202104 501362
rect 202052 501298 202104 501304
rect 202156 500818 202184 700402
rect 267660 700398 267688 703520
rect 202236 700392 202288 700398
rect 202236 700334 202288 700340
rect 267648 700392 267700 700398
rect 267648 700334 267700 700340
rect 202248 501022 202276 700334
rect 283852 700330 283880 703520
rect 300136 700777 300164 703520
rect 300122 700768 300178 700777
rect 300122 700703 300178 700712
rect 332520 700641 332548 703520
rect 332506 700632 332562 700641
rect 332506 700567 332562 700576
rect 348804 700505 348832 703520
rect 348790 700496 348846 700505
rect 348790 700431 348846 700440
rect 364996 700369 365024 703520
rect 391204 700596 391256 700602
rect 391204 700538 391256 700544
rect 364982 700360 365038 700369
rect 283840 700324 283892 700330
rect 364982 700295 365038 700304
rect 389824 700324 389876 700330
rect 283840 700266 283892 700272
rect 389824 700266 389876 700272
rect 382924 696992 382976 696998
rect 382924 696934 382976 696940
rect 291106 682816 291162 682825
rect 291106 682751 291162 682760
rect 238482 682680 238538 682689
rect 221740 682644 221792 682650
rect 238482 682615 238538 682624
rect 221740 682586 221792 682592
rect 212172 681964 212224 681970
rect 212172 681906 212224 681912
rect 207388 681760 207440 681766
rect 207388 681702 207440 681708
rect 207400 679932 207428 681702
rect 212184 679932 212212 681906
rect 216956 681896 217008 681902
rect 216956 681838 217008 681844
rect 216968 679932 216996 681838
rect 219348 681828 219400 681834
rect 219348 681770 219400 681776
rect 219360 679932 219388 681770
rect 221752 679932 221780 682586
rect 226524 682304 226576 682310
rect 226524 682246 226576 682252
rect 226536 679932 226564 682246
rect 231308 682236 231360 682242
rect 231308 682178 231360 682184
rect 231320 679932 231348 682178
rect 236092 682168 236144 682174
rect 236092 682110 236144 682116
rect 233700 682100 233752 682106
rect 233700 682042 233752 682048
rect 233712 679932 233740 682042
rect 236104 679932 236132 682110
rect 238496 679932 238524 682615
rect 255228 682576 255280 682582
rect 255228 682518 255280 682524
rect 271970 682544 272026 682553
rect 252836 682032 252888 682038
rect 252836 681974 252888 681980
rect 252848 679932 252876 681974
rect 255240 679932 255268 682518
rect 271970 682479 272026 682488
rect 276756 682508 276808 682514
rect 257620 680944 257672 680950
rect 257620 680886 257672 680892
rect 257632 679932 257660 680886
rect 262404 680876 262456 680882
rect 262404 680818 262456 680824
rect 262416 679932 262444 680818
rect 267188 680808 267240 680814
rect 267188 680750 267240 680756
rect 267200 679932 267228 680750
rect 271984 679932 272012 682479
rect 276756 682450 276808 682456
rect 274362 682408 274418 682417
rect 274362 682343 274418 682352
rect 274376 679932 274404 682343
rect 276768 679932 276796 682450
rect 279148 682440 279200 682446
rect 279148 682382 279200 682388
rect 279160 679932 279188 682382
rect 281540 682372 281592 682378
rect 281540 682314 281592 682320
rect 281552 679932 281580 682314
rect 286322 682272 286378 682281
rect 286322 682207 286378 682216
rect 283930 682136 283986 682145
rect 283930 682071 283986 682080
rect 283944 679932 283972 682071
rect 286336 679932 286364 682207
rect 288714 682000 288770 682009
rect 288714 681935 288770 681944
rect 288728 679932 288756 681935
rect 291120 679932 291148 682751
rect 317420 682712 317472 682718
rect 377772 682712 377824 682718
rect 317420 682654 317472 682660
rect 326986 682680 327042 682689
rect 303068 680740 303120 680746
rect 303068 680682 303120 680688
rect 303080 679932 303108 680682
rect 307852 680672 307904 680678
rect 307852 680614 307904 680620
rect 305458 680504 305514 680513
rect 305458 680439 305514 680448
rect 305472 679932 305500 680439
rect 307864 679932 307892 680614
rect 310244 680604 310296 680610
rect 310244 680546 310296 680552
rect 310256 679932 310284 680546
rect 312636 680536 312688 680542
rect 312636 680478 312688 680484
rect 312648 679932 312676 680478
rect 315028 680468 315080 680474
rect 315028 680410 315080 680416
rect 315040 679932 315068 680410
rect 317432 679932 317460 682654
rect 377772 682654 377824 682660
rect 326986 682615 327042 682624
rect 334164 682644 334216 682650
rect 319810 682544 319866 682553
rect 319810 682479 319866 682488
rect 322204 682508 322256 682514
rect 319824 679932 319852 682479
rect 322204 682450 322256 682456
rect 322216 679932 322244 682450
rect 327000 679932 327028 682615
rect 334164 682586 334216 682592
rect 329380 680400 329432 680406
rect 329380 680342 329432 680348
rect 331770 680368 331826 680377
rect 329392 679932 329420 680342
rect 331770 680303 331826 680312
rect 331784 679932 331812 680303
rect 334176 679932 334204 682586
rect 336556 682576 336608 682582
rect 336556 682518 336608 682524
rect 336568 679932 336596 682518
rect 355692 682440 355744 682446
rect 355692 682382 355744 682388
rect 367650 682408 367706 682417
rect 353300 682304 353352 682310
rect 341338 682272 341394 682281
rect 353300 682246 353352 682252
rect 341338 682207 341394 682216
rect 350908 682236 350960 682242
rect 338946 682136 339002 682145
rect 338946 682071 339002 682080
rect 338960 679932 338988 682071
rect 341352 679932 341380 682207
rect 350908 682178 350960 682184
rect 348516 682168 348568 682174
rect 348516 682110 348568 682116
rect 343732 682100 343784 682106
rect 343732 682042 343784 682048
rect 343744 679932 343772 682042
rect 346124 682032 346176 682038
rect 346124 681974 346176 681980
rect 346136 679932 346164 681974
rect 348528 679932 348556 682110
rect 350920 679932 350948 682178
rect 353312 679932 353340 682246
rect 355704 679932 355732 682382
rect 362868 682372 362920 682378
rect 367650 682343 367706 682352
rect 362868 682314 362920 682320
rect 360476 681896 360528 681902
rect 360476 681838 360528 681844
rect 358084 681828 358136 681834
rect 358084 681770 358136 681776
rect 358096 679932 358124 681770
rect 360488 679932 360516 681838
rect 362880 679932 362908 682314
rect 365260 681964 365312 681970
rect 365260 681906 365312 681912
rect 365272 679932 365300 681906
rect 367664 679932 367692 682343
rect 374826 682136 374882 682145
rect 374826 682071 374882 682080
rect 377588 682100 377640 682106
rect 372434 682000 372490 682009
rect 372434 681935 372490 681944
rect 370042 681864 370098 681873
rect 370042 681799 370098 681808
rect 370056 679932 370084 681799
rect 372448 679932 372476 681935
rect 374840 679932 374868 682071
rect 377588 682042 377640 682048
rect 377220 681760 377272 681766
rect 377220 681702 377272 681708
rect 377232 679932 377260 681702
rect 210976 679856 211028 679862
rect 209778 679824 209834 679833
rect 202512 679788 202564 679794
rect 202512 679730 202564 679736
rect 206008 679788 206060 679794
rect 210976 679798 211028 679804
rect 209778 679759 209834 679768
rect 206008 679730 206060 679736
rect 202524 679386 202552 679730
rect 204994 679552 205050 679561
rect 204994 679487 205050 679496
rect 206020 679454 206048 679730
rect 210988 679538 211016 679798
rect 264518 679688 264574 679697
rect 269302 679688 269358 679697
rect 264574 679646 264822 679674
rect 264518 679623 264574 679632
rect 269358 679646 269606 679674
rect 269302 679623 269358 679632
rect 259644 679584 259696 679590
rect 210988 679522 211154 679538
rect 214208 679522 214590 679538
rect 223776 679522 224158 679538
rect 247696 679522 248078 679538
rect 300674 679552 300730 679561
rect 259696 679532 260038 679538
rect 259644 679526 260038 679532
rect 210988 679516 211166 679522
rect 210988 679510 211114 679516
rect 211114 679458 211166 679464
rect 214196 679516 214590 679522
rect 214248 679510 214590 679516
rect 223764 679516 224158 679522
rect 214196 679458 214248 679464
rect 223816 679510 224158 679516
rect 247684 679516 248078 679522
rect 223764 679458 223816 679464
rect 247736 679510 248078 679516
rect 259656 679510 260038 679526
rect 300674 679487 300730 679496
rect 247684 679458 247736 679464
rect 205640 679448 205692 679454
rect 205824 679448 205876 679454
rect 205692 679396 205824 679402
rect 205640 679390 205876 679396
rect 206008 679448 206060 679454
rect 206008 679390 206060 679396
rect 228548 679448 228600 679454
rect 240508 679448 240560 679454
rect 228600 679396 228942 679402
rect 228548 679390 228942 679396
rect 242900 679448 242952 679454
rect 240560 679396 240902 679402
rect 240508 679390 240902 679396
rect 245568 679448 245620 679454
rect 242952 679396 243294 679402
rect 242900 679390 243294 679396
rect 250076 679448 250128 679454
rect 245620 679396 245686 679402
rect 245568 679390 245686 679396
rect 324872 679448 324924 679454
rect 293498 679416 293554 679425
rect 250128 679396 250470 679402
rect 250076 679390 250470 679396
rect 202512 679380 202564 679386
rect 205652 679374 205864 679390
rect 228560 679374 228942 679390
rect 240520 679374 240902 679390
rect 242912 679374 243294 679390
rect 245580 679374 245686 679390
rect 250088 679374 250470 679390
rect 324622 679396 324872 679402
rect 324622 679390 324924 679396
rect 324622 679374 324912 679390
rect 293498 679351 293554 679360
rect 202512 679322 202564 679328
rect 295890 679280 295946 679289
rect 202340 679250 202630 679266
rect 202328 679244 202630 679250
rect 202380 679238 202630 679244
rect 295890 679215 295946 679224
rect 298282 679280 298338 679289
rect 298282 679215 298338 679224
rect 202328 679186 202380 679192
rect 202328 678836 202380 678842
rect 202328 678778 202380 678784
rect 202236 501016 202288 501022
rect 202236 500958 202288 500964
rect 202144 500812 202196 500818
rect 202144 500754 202196 500760
rect 201960 500744 202012 500750
rect 201960 500686 202012 500692
rect 201592 496256 201644 496262
rect 201592 496198 201644 496204
rect 201500 481092 201552 481098
rect 201500 481034 201552 481040
rect 202340 466070 202368 678778
rect 202420 678360 202472 678366
rect 202420 678302 202472 678308
rect 202432 466342 202460 678302
rect 207572 500744 207624 500750
rect 203076 500670 203196 500698
rect 207572 500686 207624 500692
rect 213368 500744 213420 500750
rect 214288 500744 214340 500750
rect 213368 500686 213420 500692
rect 213918 500712 213974 500721
rect 203076 500614 203104 500670
rect 203168 500614 203196 500670
rect 203064 500608 203116 500614
rect 203064 500550 203116 500556
rect 203156 500608 203208 500614
rect 203156 500550 203208 500556
rect 203156 500472 203208 500478
rect 203340 500472 203392 500478
rect 203208 500420 203340 500426
rect 203156 500414 203392 500420
rect 203168 500398 203380 500414
rect 207584 500138 207612 500686
rect 212538 500304 212594 500313
rect 212538 500239 212594 500248
rect 211158 500168 211214 500177
rect 207572 500132 207624 500138
rect 211158 500103 211214 500112
rect 207572 500074 207624 500080
rect 207020 498908 207072 498914
rect 207020 498850 207072 498856
rect 205640 483676 205692 483682
rect 205640 483618 205692 483624
rect 204260 470620 204312 470626
rect 204260 470562 204312 470568
rect 202420 466336 202472 466342
rect 202420 466278 202472 466284
rect 202328 466064 202380 466070
rect 202328 466006 202380 466012
rect 201408 465656 201460 465662
rect 201408 465598 201460 465604
rect 201040 463140 201092 463146
rect 201040 463082 201092 463088
rect 200856 461780 200908 461786
rect 200856 461722 200908 461728
rect 204272 460934 204300 470562
rect 200776 460906 200896 460934
rect 204272 460906 205220 460934
rect 200028 460692 200080 460698
rect 200028 460634 200080 460640
rect 200672 456476 200724 456482
rect 200672 456418 200724 456424
rect 200304 454504 200356 454510
rect 200304 454446 200356 454452
rect 199304 449942 199594 449970
rect 199672 449942 199962 449970
rect 200316 449956 200344 454446
rect 200684 449956 200712 456418
rect 200868 453626 200896 460906
rect 201500 457360 201552 457366
rect 201500 457302 201552 457308
rect 201512 456794 201540 457302
rect 204352 456952 204404 456958
rect 204352 456894 204404 456900
rect 203064 456884 203116 456890
rect 203064 456826 203116 456832
rect 201512 456766 201908 456794
rect 201776 455592 201828 455598
rect 201776 455534 201828 455540
rect 201040 455524 201092 455530
rect 201040 455466 201092 455472
rect 200856 453620 200908 453626
rect 200856 453562 200908 453568
rect 201052 449956 201080 455466
rect 201406 451480 201462 451489
rect 201406 451415 201462 451424
rect 201420 449956 201448 451415
rect 201788 449956 201816 455534
rect 201880 449970 201908 456766
rect 202512 455660 202564 455666
rect 202512 455602 202564 455608
rect 201880 449942 202170 449970
rect 202524 449956 202552 455602
rect 202880 454572 202932 454578
rect 202880 454514 202932 454520
rect 202892 449956 202920 454514
rect 203076 449970 203104 456826
rect 203616 452328 203668 452334
rect 203616 452270 203668 452276
rect 203076 449942 203274 449970
rect 203628 449956 203656 452270
rect 203984 452260 204036 452266
rect 203984 452202 204036 452208
rect 203996 449956 204024 452202
rect 204260 451240 204312 451246
rect 204260 451182 204312 451188
rect 204272 450566 204300 451182
rect 204260 450560 204312 450566
rect 204260 450502 204312 450508
rect 204364 449956 204392 456894
rect 204812 456816 204864 456822
rect 204812 456758 204864 456764
rect 204720 455728 204772 455734
rect 204720 455670 204772 455676
rect 204732 449956 204760 455670
rect 204824 449970 204852 456758
rect 205192 449970 205220 460906
rect 205652 456074 205680 483618
rect 205732 482316 205784 482322
rect 205732 482258 205784 482264
rect 205640 456068 205692 456074
rect 205640 456010 205692 456016
rect 205744 455682 205772 482258
rect 205824 478168 205876 478174
rect 205824 478110 205876 478116
rect 205836 455938 205864 478110
rect 205916 474020 205968 474026
rect 205916 473962 205968 473968
rect 205928 460934 205956 473962
rect 205928 460906 206140 460934
rect 205824 455932 205876 455938
rect 205824 455874 205876 455880
rect 205744 455654 206048 455682
rect 205916 451308 205968 451314
rect 205916 451250 205968 451256
rect 205928 449970 205956 451250
rect 204824 449942 205114 449970
rect 205192 449942 205482 449970
rect 205850 449942 205956 449970
rect 206020 449970 206048 455654
rect 206112 451314 206140 460906
rect 206284 456068 206336 456074
rect 206284 456010 206336 456016
rect 206100 451308 206152 451314
rect 206100 451250 206152 451256
rect 206296 449970 206324 456010
rect 206652 455932 206704 455938
rect 206652 455874 206704 455880
rect 206664 449970 206692 455874
rect 207032 449970 207060 498850
rect 207112 494760 207164 494766
rect 207112 494702 207164 494708
rect 207124 460934 207152 494702
rect 208400 493332 208452 493338
rect 208400 493274 208452 493280
rect 207124 460906 207428 460934
rect 207400 449970 207428 460906
rect 207756 457496 207808 457502
rect 207756 457438 207808 457444
rect 207768 449970 207796 457438
rect 206020 449942 206218 449970
rect 206296 449942 206586 449970
rect 206664 449942 206954 449970
rect 207032 449942 207322 449970
rect 207400 449942 207690 449970
rect 207768 449942 208058 449970
rect 208412 449956 208440 493274
rect 208492 492108 208544 492114
rect 208492 492050 208544 492056
rect 208504 456074 208532 492050
rect 209780 490816 209832 490822
rect 209780 490758 209832 490764
rect 208584 486464 208636 486470
rect 208584 486406 208636 486412
rect 208492 456068 208544 456074
rect 208492 456010 208544 456016
rect 208596 449970 208624 486406
rect 209044 484424 209096 484430
rect 209044 484366 209096 484372
rect 208860 457564 208912 457570
rect 208860 457506 208912 457512
rect 208872 449970 208900 457506
rect 209056 456822 209084 484366
rect 209136 457360 209188 457366
rect 209136 457302 209188 457308
rect 209148 456822 209176 457302
rect 209044 456816 209096 456822
rect 209044 456758 209096 456764
rect 209136 456816 209188 456822
rect 209136 456758 209188 456764
rect 209504 456476 209556 456482
rect 209504 456418 209556 456424
rect 209228 456068 209280 456074
rect 209228 456010 209280 456016
rect 209320 456068 209372 456074
rect 209320 456010 209372 456016
rect 209240 449970 209268 456010
rect 209332 455734 209360 456010
rect 209320 455728 209372 455734
rect 209320 455670 209372 455676
rect 209412 455728 209464 455734
rect 209412 455670 209464 455676
rect 209424 455598 209452 455670
rect 209516 455598 209544 456418
rect 209412 455592 209464 455598
rect 209412 455534 209464 455540
rect 209504 455592 209556 455598
rect 209504 455534 209556 455540
rect 209792 449970 209820 490758
rect 209870 480856 209926 480865
rect 209870 480791 209926 480800
rect 209884 455938 209912 480791
rect 209964 475584 210016 475590
rect 209964 475526 210016 475532
rect 209976 460934 210004 475526
rect 209976 460906 210372 460934
rect 210056 457768 210108 457774
rect 210056 457710 210108 457716
rect 209872 455932 209924 455938
rect 209872 455874 209924 455880
rect 210068 449970 210096 457710
rect 210344 449970 210372 460906
rect 210700 455932 210752 455938
rect 210700 455874 210752 455880
rect 210712 449970 210740 455874
rect 211172 449970 211200 500103
rect 211250 497448 211306 497457
rect 211250 497383 211306 497392
rect 211264 455938 211292 497383
rect 211342 462904 211398 462913
rect 211342 462839 211398 462848
rect 211356 460934 211384 462839
rect 211356 460906 211844 460934
rect 211434 457464 211490 457473
rect 211434 457399 211490 457408
rect 211252 455932 211304 455938
rect 211252 455874 211304 455880
rect 211448 449970 211476 457399
rect 211816 449970 211844 460906
rect 212172 455932 212224 455938
rect 212172 455874 212224 455880
rect 212184 449970 212212 455874
rect 212552 450158 212580 500239
rect 213380 500206 213408 500686
rect 213918 500647 213974 500656
rect 214102 500712 214158 500721
rect 215576 500744 215628 500750
rect 214288 500686 214340 500692
rect 215404 500692 215576 500698
rect 215404 500686 215628 500692
rect 215668 500744 215720 500750
rect 215668 500686 215720 500692
rect 228364 500744 228416 500750
rect 228364 500686 228416 500692
rect 349344 500744 349396 500750
rect 349344 500686 349396 500692
rect 351828 500744 351880 500750
rect 354864 500744 354916 500750
rect 351828 500686 351880 500692
rect 354862 500712 354864 500721
rect 354956 500744 355008 500750
rect 354916 500712 354918 500721
rect 214102 500647 214158 500656
rect 213368 500200 213420 500206
rect 213368 500142 213420 500148
rect 212630 499896 212686 499905
rect 212630 499831 212686 499840
rect 212540 450152 212592 450158
rect 212540 450094 212592 450100
rect 212644 450090 212672 499831
rect 212724 496188 212776 496194
rect 212724 496130 212776 496136
rect 212632 450084 212684 450090
rect 212632 450026 212684 450032
rect 212736 449970 212764 496130
rect 212908 450152 212960 450158
rect 212908 450094 212960 450100
rect 212920 449970 212948 450094
rect 213276 450084 213328 450090
rect 213276 450026 213328 450032
rect 213288 449970 213316 450026
rect 208596 449942 208794 449970
rect 208872 449942 209162 449970
rect 209240 449942 209530 449970
rect 209792 449942 209898 449970
rect 210068 449942 210266 449970
rect 210344 449942 210634 449970
rect 210712 449942 211002 449970
rect 211172 449942 211370 449970
rect 211448 449942 211738 449970
rect 211816 449942 212106 449970
rect 212184 449942 212474 449970
rect 212736 449942 212842 449970
rect 212920 449942 213210 449970
rect 213288 449942 213578 449970
rect 213932 449956 213960 500647
rect 214010 500576 214066 500585
rect 214010 500511 214066 500520
rect 214024 449970 214052 500511
rect 214116 450106 214144 500647
rect 214300 492674 214328 500686
rect 215404 500670 215616 500686
rect 215298 500032 215354 500041
rect 215298 499967 215354 499976
rect 214208 492646 214328 492674
rect 214208 460934 214236 492646
rect 214208 460906 214788 460934
rect 214564 452328 214616 452334
rect 214564 452270 214616 452276
rect 214472 452260 214524 452266
rect 214472 452202 214524 452208
rect 214484 451586 214512 452202
rect 214576 451654 214604 452270
rect 214564 451648 214616 451654
rect 214564 451590 214616 451596
rect 214472 451580 214524 451586
rect 214472 451522 214524 451528
rect 214116 450078 214420 450106
rect 214392 449970 214420 450078
rect 214760 449970 214788 460906
rect 215312 450158 215340 499967
rect 215300 450152 215352 450158
rect 215300 450094 215352 450100
rect 214024 449942 214314 449970
rect 214392 449942 214682 449970
rect 214760 449942 215050 449970
rect 215404 449956 215432 500670
rect 215484 500200 215536 500206
rect 215484 500142 215536 500148
rect 215496 449970 215524 500142
rect 215680 500138 215708 500686
rect 216956 500676 217008 500682
rect 216956 500618 217008 500624
rect 215668 500132 215720 500138
rect 215668 500074 215720 500080
rect 215576 481092 215628 481098
rect 215576 481034 215628 481040
rect 215588 460934 215616 481034
rect 216772 461916 216824 461922
rect 216772 461858 216824 461864
rect 215588 460906 215892 460934
rect 215864 449970 215892 460906
rect 216680 459060 216732 459066
rect 216680 459002 216732 459008
rect 216692 450158 216720 459002
rect 216220 450152 216272 450158
rect 216220 450094 216272 450100
rect 216680 450152 216732 450158
rect 216680 450094 216732 450100
rect 216232 449970 216260 450094
rect 216784 450090 216812 461858
rect 216864 461848 216916 461854
rect 216864 461790 216916 461796
rect 216772 450084 216824 450090
rect 216772 450026 216824 450032
rect 215496 449942 215786 449970
rect 215864 449942 216154 449970
rect 216232 449942 216522 449970
rect 216876 449956 216904 461790
rect 216968 449970 216996 500618
rect 219440 500540 219492 500546
rect 219440 500482 219492 500488
rect 218058 468480 218114 468489
rect 218058 468415 218114 468424
rect 218072 462482 218100 468415
rect 217980 462454 218100 462482
rect 217980 461700 218008 462454
rect 218060 462392 218112 462398
rect 218060 462334 218112 462340
rect 218072 461854 218100 462334
rect 218152 461984 218204 461990
rect 218152 461926 218204 461932
rect 218060 461848 218112 461854
rect 218060 461790 218112 461796
rect 217980 461672 218100 461700
rect 217324 450152 217376 450158
rect 217324 450094 217376 450100
rect 217336 449970 217364 450094
rect 217692 450084 217744 450090
rect 217692 450026 217744 450032
rect 217704 449970 217732 450026
rect 218072 449970 218100 461672
rect 218164 450158 218192 461926
rect 218428 459128 218480 459134
rect 218428 459070 218480 459076
rect 218152 450152 218204 450158
rect 218152 450094 218204 450100
rect 218440 449970 218468 459070
rect 219452 450566 219480 500482
rect 219532 498976 219584 498982
rect 219532 498918 219584 498924
rect 219440 450560 219492 450566
rect 219440 450502 219492 450508
rect 219544 450158 219572 498918
rect 221096 485172 221148 485178
rect 221096 485114 221148 485120
rect 220912 475516 220964 475522
rect 220912 475458 220964 475464
rect 219624 471436 219676 471442
rect 219624 471378 219676 471384
rect 219636 451042 219664 471378
rect 219716 461712 219768 461718
rect 219716 461654 219768 461660
rect 219624 451036 219676 451042
rect 219624 450978 219676 450984
rect 218796 450152 218848 450158
rect 218796 450094 218848 450100
rect 219532 450152 219584 450158
rect 219532 450094 219584 450100
rect 218808 449970 218836 450094
rect 216968 449942 217258 449970
rect 217336 449942 217626 449970
rect 217704 449942 217994 449970
rect 218072 449942 218362 449970
rect 218440 449942 218730 449970
rect 218808 449942 219098 449970
rect 193864 449880 193916 449886
rect 219728 449834 219756 461654
rect 220820 457632 220872 457638
rect 220820 457574 220872 457580
rect 219808 451036 219860 451042
rect 219808 450978 219860 450984
rect 219820 449956 219848 450978
rect 219900 450560 219952 450566
rect 219900 450502 219952 450508
rect 219912 449970 219940 450502
rect 220268 450152 220320 450158
rect 220268 450094 220320 450100
rect 220280 449970 220308 450094
rect 220832 450090 220860 457574
rect 220924 450566 220952 475458
rect 221004 457700 221056 457706
rect 221004 457642 221056 457648
rect 220912 450560 220964 450566
rect 220912 450502 220964 450508
rect 221016 450158 221044 457642
rect 221004 450152 221056 450158
rect 221004 450094 221056 450100
rect 220820 450084 220872 450090
rect 220820 450026 220872 450032
rect 221108 449970 221136 485114
rect 222476 483812 222528 483818
rect 222476 483754 222528 483760
rect 222292 461644 222344 461650
rect 222292 461586 222344 461592
rect 222200 456136 222252 456142
rect 222200 456078 222252 456084
rect 221372 450560 221424 450566
rect 221372 450502 221424 450508
rect 221188 450084 221240 450090
rect 221188 450026 221240 450032
rect 219912 449942 220202 449970
rect 220280 449942 220570 449970
rect 220938 449942 221136 449970
rect 221200 449970 221228 450026
rect 221384 449970 221412 450502
rect 222212 450158 222240 456078
rect 221740 450152 221792 450158
rect 221740 450094 221792 450100
rect 222200 450152 222252 450158
rect 222200 450094 222252 450100
rect 221752 449970 221780 450094
rect 222304 449970 222332 461586
rect 222488 460934 222516 483754
rect 225052 461848 225104 461854
rect 225052 461790 225104 461796
rect 222488 460906 222884 460934
rect 222476 458856 222528 458862
rect 222476 458798 222528 458804
rect 222488 449970 222516 458798
rect 222856 449970 222884 460906
rect 223948 460216 224000 460222
rect 223948 460158 224000 460164
rect 223672 458924 223724 458930
rect 223672 458866 223724 458872
rect 223212 450152 223264 450158
rect 223212 450094 223264 450100
rect 223224 449970 223252 450094
rect 223684 449970 223712 458866
rect 223960 449970 223988 460158
rect 224316 457836 224368 457842
rect 224316 457778 224368 457784
rect 224328 449970 224356 457778
rect 224960 453212 225012 453218
rect 224960 453154 225012 453160
rect 221200 449942 221306 449970
rect 221384 449942 221674 449970
rect 221752 449942 222042 449970
rect 222304 449942 222410 449970
rect 222488 449942 222778 449970
rect 222856 449942 223146 449970
rect 223224 449942 223514 449970
rect 223684 449942 223882 449970
rect 223960 449942 224250 449970
rect 224328 449942 224618 449970
rect 224972 449956 225000 453154
rect 225064 449970 225092 461790
rect 227996 454980 228048 454986
rect 227996 454922 228048 454928
rect 227260 454912 227312 454918
rect 227260 454854 227312 454860
rect 226800 452124 226852 452130
rect 226800 452066 226852 452072
rect 226432 451308 226484 451314
rect 226432 451250 226484 451256
rect 226064 450764 226116 450770
rect 226064 450706 226116 450712
rect 225064 449942 225354 449970
rect 225524 449954 225722 449970
rect 226076 449956 226104 450706
rect 226444 449956 226472 451250
rect 226812 449956 226840 452066
rect 227168 451852 227220 451858
rect 227168 451794 227220 451800
rect 227180 449956 227208 451794
rect 227272 449970 227300 454854
rect 227904 450696 227956 450702
rect 227904 450638 227956 450644
rect 225512 449948 225722 449954
rect 225564 449942 225722 449948
rect 227272 449942 227562 449970
rect 227916 449956 227944 450638
rect 228008 449970 228036 454922
rect 228376 452538 228404 500686
rect 346400 500676 346452 500682
rect 346400 500618 346452 500624
rect 238760 500608 238812 500614
rect 343640 500608 343692 500614
rect 238760 500550 238812 500556
rect 320178 500576 320234 500585
rect 228454 500440 228510 500449
rect 228454 500375 228510 500384
rect 228364 452532 228416 452538
rect 228364 452474 228416 452480
rect 228468 452470 228496 500375
rect 228548 498160 228600 498166
rect 228548 498102 228600 498108
rect 237654 498128 237710 498137
rect 228456 452464 228508 452470
rect 228456 452406 228508 452412
rect 228560 452266 228588 498102
rect 228640 498092 228692 498098
rect 237654 498063 237710 498072
rect 228640 498034 228692 498040
rect 228548 452260 228600 452266
rect 228548 452202 228600 452208
rect 228652 452062 228680 498034
rect 234710 497584 234766 497593
rect 234710 497519 234766 497528
rect 228732 497412 228784 497418
rect 228732 497354 228784 497360
rect 228744 452402 228772 497354
rect 232504 495032 232556 495038
rect 232504 494974 232556 494980
rect 231308 454232 231360 454238
rect 231308 454174 231360 454180
rect 230110 453384 230166 453393
rect 230110 453319 230166 453328
rect 229744 453144 229796 453150
rect 229744 453086 229796 453092
rect 229376 453076 229428 453082
rect 229376 453018 229428 453024
rect 228732 452396 228784 452402
rect 228732 452338 228784 452344
rect 228364 452056 228416 452062
rect 228364 451998 228416 452004
rect 228640 452056 228692 452062
rect 228640 451998 228692 452004
rect 228376 449970 228404 451998
rect 228916 451988 228968 451994
rect 228916 451930 228968 451936
rect 228928 451274 228956 451930
rect 228928 451246 229048 451274
rect 228008 449942 228298 449970
rect 228376 449942 228666 449970
rect 229020 449956 229048 451246
rect 229388 449956 229416 453018
rect 229756 449956 229784 453086
rect 230124 449956 230152 453319
rect 231216 451376 231268 451382
rect 231216 451318 231268 451324
rect 230848 450628 230900 450634
rect 230848 450570 230900 450576
rect 230860 449956 230888 450570
rect 231228 449956 231256 451318
rect 231320 449970 231348 454174
rect 232516 451926 232544 494974
rect 232596 494964 232648 494970
rect 232596 494906 232648 494912
rect 232608 452334 232636 494906
rect 232688 464500 232740 464506
rect 232688 464442 232740 464448
rect 232596 452328 232648 452334
rect 232596 452270 232648 452276
rect 232700 452130 232728 464442
rect 232780 464432 232832 464438
rect 232780 464374 232832 464380
rect 232792 460934 232820 464374
rect 234724 460934 234752 497519
rect 235264 496256 235316 496262
rect 235264 496198 235316 496204
rect 232792 460906 232912 460934
rect 234724 460906 235212 460934
rect 232778 454336 232834 454345
rect 232778 454271 232834 454280
rect 232688 452124 232740 452130
rect 232688 452066 232740 452072
rect 231952 451920 232004 451926
rect 231952 451862 232004 451868
rect 232504 451920 232556 451926
rect 232504 451862 232556 451868
rect 231320 449942 231610 449970
rect 231964 449956 231992 451862
rect 232688 451716 232740 451722
rect 232688 451658 232740 451664
rect 232320 451512 232372 451518
rect 232320 451454 232372 451460
rect 232332 449956 232360 451454
rect 232700 449956 232728 451658
rect 232792 449970 232820 454271
rect 232884 452062 232912 460906
rect 233884 454300 233936 454306
rect 233884 454242 233936 454248
rect 233516 454164 233568 454170
rect 233516 454106 233568 454112
rect 232872 452056 232924 452062
rect 232872 451998 232924 452004
rect 233422 449984 233478 449993
rect 232792 449942 233082 449970
rect 233528 449970 233556 454106
rect 233896 449970 233924 454242
rect 234894 452296 234950 452305
rect 234894 452231 234950 452240
rect 234528 451444 234580 451450
rect 234528 451386 234580 451392
rect 233528 449942 233818 449970
rect 233896 449942 234186 449970
rect 234540 449956 234568 451386
rect 234908 449956 234936 452231
rect 234988 452192 235040 452198
rect 234988 452134 235040 452140
rect 235000 449970 235028 452134
rect 235184 450106 235212 460906
rect 235276 452606 235304 496198
rect 237472 465588 237524 465594
rect 237472 465530 237524 465536
rect 235356 464296 235408 464302
rect 235356 464238 235408 464244
rect 235264 452600 235316 452606
rect 235264 452542 235316 452548
rect 235368 452198 235396 464238
rect 236184 462868 236236 462874
rect 236184 462810 236236 462816
rect 236196 460934 236224 462810
rect 236196 460906 236500 460934
rect 236368 452600 236420 452606
rect 236368 452542 236420 452548
rect 235356 452192 235408 452198
rect 235356 452134 235408 452140
rect 235998 452160 236054 452169
rect 235998 452095 236054 452104
rect 235184 450078 235396 450106
rect 235368 449970 235396 450078
rect 235000 449942 235290 449970
rect 235368 449942 235658 449970
rect 236012 449956 236040 452095
rect 236380 449956 236408 452542
rect 236472 449970 236500 460906
rect 237484 453082 237512 465530
rect 237472 453076 237524 453082
rect 237472 453018 237524 453024
rect 237104 452532 237156 452538
rect 237104 452474 237156 452480
rect 236472 449942 236762 449970
rect 237116 449956 237144 452474
rect 237668 449970 237696 498063
rect 237932 460692 237984 460698
rect 237932 460634 237984 460640
rect 237840 452464 237892 452470
rect 237840 452406 237892 452412
rect 237498 449942 237696 449970
rect 237852 449956 237880 452406
rect 237944 449970 237972 460634
rect 238772 453082 238800 500550
rect 343640 500550 343692 500556
rect 320178 500511 320234 500520
rect 336740 500540 336792 500546
rect 242900 500472 242952 500478
rect 242900 500414 242952 500420
rect 288438 500440 288494 500449
rect 241520 500404 241572 500410
rect 241520 500346 241572 500352
rect 238852 498024 238904 498030
rect 238852 497966 238904 497972
rect 238942 497992 238998 498001
rect 238300 453076 238352 453082
rect 238300 453018 238352 453024
rect 238760 453076 238812 453082
rect 238760 453018 238812 453024
rect 238312 449970 238340 453018
rect 238864 449970 238892 497966
rect 238942 497927 238998 497936
rect 238956 456794 238984 497927
rect 240140 497548 240192 497554
rect 240140 497490 240192 497496
rect 240232 497548 240284 497554
rect 240232 497490 240284 497496
rect 239036 462936 239088 462942
rect 239036 462878 239088 462884
rect 239048 460934 239076 462878
rect 239048 460906 239812 460934
rect 238956 456766 239076 456794
rect 239048 449970 239076 456766
rect 239404 453076 239456 453082
rect 239404 453018 239456 453024
rect 239416 449970 239444 453018
rect 239784 449970 239812 460906
rect 240152 453082 240180 497490
rect 240244 453150 240272 497490
rect 240324 465656 240376 465662
rect 240324 465598 240376 465604
rect 240336 460934 240364 465598
rect 240336 460906 240548 460934
rect 240232 453144 240284 453150
rect 240232 453086 240284 453092
rect 240140 453076 240192 453082
rect 240140 453018 240192 453024
rect 240520 449970 240548 460906
rect 240876 453144 240928 453150
rect 240876 453086 240928 453092
rect 240600 453076 240652 453082
rect 240600 453018 240652 453024
rect 237944 449942 238234 449970
rect 238312 449942 238602 449970
rect 238864 449942 238970 449970
rect 239048 449942 239338 449970
rect 239416 449942 239706 449970
rect 239784 449942 240074 449970
rect 240442 449942 240548 449970
rect 240612 449970 240640 453018
rect 240888 449970 240916 453086
rect 240612 449942 240810 449970
rect 240888 449942 241178 449970
rect 241532 449956 241560 500346
rect 241612 497616 241664 497622
rect 241612 497558 241664 497564
rect 241624 453150 241652 497558
rect 241704 466404 241756 466410
rect 241704 466346 241756 466352
rect 241612 453144 241664 453150
rect 241612 453086 241664 453092
rect 241716 453082 241744 466346
rect 241796 463684 241848 463690
rect 241796 463626 241848 463632
rect 241704 453076 241756 453082
rect 241704 453018 241756 453024
rect 241808 449970 241836 463626
rect 242348 453144 242400 453150
rect 242348 453086 242400 453092
rect 241980 453076 242032 453082
rect 241980 453018 242032 453024
rect 241992 449970 242020 453018
rect 242360 449970 242388 453086
rect 242912 451110 242940 500414
rect 288438 500375 288494 500384
rect 244280 500336 244332 500342
rect 244280 500278 244332 500284
rect 242992 497616 243044 497622
rect 242992 497558 243044 497564
rect 242900 451104 242952 451110
rect 242900 451046 242952 451052
rect 243004 450922 243032 497558
rect 243084 466268 243136 466274
rect 243084 466210 243136 466216
rect 243096 453082 243124 466210
rect 243176 463616 243228 463622
rect 243176 463558 243228 463564
rect 243188 460934 243216 463558
rect 243188 460906 243492 460934
rect 243084 453076 243136 453082
rect 243084 453018 243136 453024
rect 243360 451104 243412 451110
rect 243360 451046 243412 451052
rect 243004 450894 243124 450922
rect 243096 449970 243124 450894
rect 241808 449942 241914 449970
rect 241992 449942 242282 449970
rect 242360 449942 242650 449970
rect 243018 449942 243124 449970
rect 243372 449956 243400 451046
rect 243464 449970 243492 460906
rect 244292 453082 244320 500278
rect 254216 500268 254268 500274
rect 254216 500210 254268 500216
rect 244936 499526 244964 500140
rect 244924 499520 244976 499526
rect 244922 499488 244924 499497
rect 244976 499488 244978 499497
rect 244922 499423 244978 499432
rect 244936 499397 244964 499423
rect 249800 499112 249852 499118
rect 249800 499054 249852 499060
rect 247038 497856 247094 497865
rect 247038 497791 247094 497800
rect 245658 497720 245714 497729
rect 244372 497684 244424 497690
rect 245658 497655 245714 497664
rect 244372 497626 244424 497632
rect 243820 453076 243872 453082
rect 243820 453018 243872 453024
rect 244280 453076 244332 453082
rect 244280 453018 244332 453024
rect 243832 449970 243860 453018
rect 244384 449970 244412 497626
rect 244462 494864 244518 494873
rect 244462 494799 244518 494808
rect 244476 456794 244504 494799
rect 244556 463548 244608 463554
rect 244556 463490 244608 463496
rect 244568 460934 244596 463490
rect 244568 460906 245332 460934
rect 244476 456766 244596 456794
rect 244568 449970 244596 456766
rect 244924 453076 244976 453082
rect 244924 453018 244976 453024
rect 244936 449970 244964 453018
rect 245304 449970 245332 460906
rect 245672 453082 245700 497655
rect 245750 494728 245806 494737
rect 245750 494663 245806 494672
rect 245764 453150 245792 494663
rect 245844 466132 245896 466138
rect 245844 466074 245896 466080
rect 245856 460934 245884 466074
rect 245856 460906 246068 460934
rect 245752 453144 245804 453150
rect 245752 453086 245804 453092
rect 245660 453076 245712 453082
rect 245660 453018 245712 453024
rect 246040 449970 246068 460906
rect 247052 453150 247080 497791
rect 247132 497752 247184 497758
rect 247132 497694 247184 497700
rect 246396 453144 246448 453150
rect 246396 453086 246448 453092
rect 247040 453144 247092 453150
rect 247040 453086 247092 453092
rect 246120 453076 246172 453082
rect 246120 453018 246172 453024
rect 243464 449942 243754 449970
rect 243832 449942 244122 449970
rect 244384 449942 244490 449970
rect 244568 449942 244858 449970
rect 244936 449942 245226 449970
rect 245304 449942 245594 449970
rect 245962 449942 246068 449970
rect 246132 449970 246160 453018
rect 246408 449970 246436 453086
rect 247144 449970 247172 497694
rect 248420 495100 248472 495106
rect 248420 495042 248472 495048
rect 247224 466200 247276 466206
rect 247224 466142 247276 466148
rect 247236 453082 247264 466142
rect 247316 463480 247368 463486
rect 247316 463422 247368 463428
rect 247224 453076 247276 453082
rect 247224 453018 247276 453024
rect 246132 449942 246330 449970
rect 246408 449942 246698 449970
rect 247066 449942 247172 449970
rect 247328 449970 247356 463422
rect 247868 453144 247920 453150
rect 247868 453086 247920 453092
rect 247500 453076 247552 453082
rect 247500 453018 247552 453024
rect 247512 449970 247540 453018
rect 247880 449970 247908 453086
rect 248432 449970 248460 495042
rect 248512 466336 248564 466342
rect 248512 466278 248564 466284
rect 248524 458266 248552 466278
rect 248602 466168 248658 466177
rect 248602 466103 248658 466112
rect 248616 460934 248644 466103
rect 248616 460906 249380 460934
rect 248524 458238 249012 458266
rect 248878 452568 248934 452577
rect 248878 452503 248934 452512
rect 247328 449942 247434 449970
rect 247512 449942 247802 449970
rect 247880 449942 248170 449970
rect 248432 449942 248538 449970
rect 248892 449956 248920 452503
rect 248984 449970 249012 458238
rect 249352 449970 249380 460906
rect 249812 449970 249840 499054
rect 251180 499044 251232 499050
rect 251180 498986 251232 498992
rect 249892 495032 249944 495038
rect 249892 494974 249944 494980
rect 249904 450106 249932 494974
rect 249984 468648 250036 468654
rect 249984 468590 250036 468596
rect 249996 453082 250024 468590
rect 250076 465928 250128 465934
rect 250076 465870 250128 465876
rect 250088 460934 250116 465870
rect 250088 460906 250484 460934
rect 249984 453076 250036 453082
rect 249984 453018 250036 453024
rect 249904 450078 250116 450106
rect 250088 449970 250116 450078
rect 250456 449970 250484 460906
rect 250812 453076 250864 453082
rect 250812 453018 250864 453024
rect 250824 449970 250852 453018
rect 251192 449970 251220 498986
rect 254032 497684 254084 497690
rect 254032 497626 254084 497632
rect 252836 495168 252888 495174
rect 252836 495110 252888 495116
rect 251272 494964 251324 494970
rect 251272 494906 251324 494912
rect 251284 456794 251312 494906
rect 252652 468716 252704 468722
rect 252652 468658 252704 468664
rect 251364 465996 251416 466002
rect 251364 465938 251416 465944
rect 251376 460934 251404 465938
rect 251376 460906 251956 460934
rect 251284 456766 251588 456794
rect 251560 449970 251588 456766
rect 251928 449970 251956 460906
rect 252664 449970 252692 468658
rect 252744 466064 252796 466070
rect 252744 466006 252796 466012
rect 252756 453082 252784 466006
rect 252848 460934 252876 495110
rect 252848 460906 253060 460934
rect 252744 453076 252796 453082
rect 252744 453018 252796 453024
rect 252928 452328 252980 452334
rect 252928 452270 252980 452276
rect 248984 449942 249274 449970
rect 249352 449942 249642 449970
rect 249812 449942 250010 449970
rect 250088 449942 250378 449970
rect 250456 449942 250746 449970
rect 250824 449942 251114 449970
rect 251192 449942 251482 449970
rect 251560 449942 251850 449970
rect 251928 449942 252218 449970
rect 252586 449942 252692 449970
rect 252940 449956 252968 452270
rect 253032 449970 253060 460906
rect 254044 456142 254072 497626
rect 254124 463412 254176 463418
rect 254124 463354 254176 463360
rect 254032 456136 254084 456142
rect 254032 456078 254084 456084
rect 253388 453076 253440 453082
rect 253388 453018 253440 453024
rect 253400 449970 253428 453018
rect 254136 449970 254164 463354
rect 254228 460934 254256 500210
rect 261024 498976 261076 498982
rect 261024 498918 261076 498924
rect 259644 498092 259696 498098
rect 259644 498034 259696 498040
rect 258172 498024 258224 498030
rect 258172 497966 258224 497972
rect 256700 497888 256752 497894
rect 256700 497830 256752 497836
rect 255412 497820 255464 497826
rect 255412 497762 255464 497768
rect 254228 460906 254900 460934
rect 254492 456136 254544 456142
rect 254492 456078 254544 456084
rect 254400 451920 254452 451926
rect 254400 451862 254452 451868
rect 253032 449942 253322 449970
rect 253400 449942 253690 449970
rect 254058 449942 254164 449970
rect 254412 449956 254440 451862
rect 254504 449970 254532 456078
rect 254872 449970 254900 460906
rect 255424 456142 255452 497762
rect 255596 497752 255648 497758
rect 255596 497694 255648 497700
rect 255608 460934 255636 497694
rect 255608 460906 256004 460934
rect 255412 456136 255464 456142
rect 255412 456078 255464 456084
rect 255504 451988 255556 451994
rect 255504 451930 255556 451936
rect 254504 449942 254794 449970
rect 254872 449942 255162 449970
rect 255516 449956 255544 451930
rect 255872 451920 255924 451926
rect 255872 451862 255924 451868
rect 255884 449956 255912 451862
rect 255976 449970 256004 460906
rect 256332 456136 256384 456142
rect 256332 456078 256384 456084
rect 256344 449970 256372 456078
rect 256712 449970 256740 497830
rect 256792 497820 256844 497826
rect 256792 497762 256844 497768
rect 256804 460934 256832 497762
rect 256804 460906 257476 460934
rect 257344 451988 257396 451994
rect 257344 451930 257396 451936
rect 255976 449942 256266 449970
rect 256344 449942 256634 449970
rect 256712 449942 257002 449970
rect 257356 449956 257384 451930
rect 257448 449970 257476 460906
rect 258184 456142 258212 497966
rect 259460 497956 259512 497962
rect 259460 497898 259512 497904
rect 259552 497956 259604 497962
rect 259552 497898 259604 497904
rect 258264 497888 258316 497894
rect 258264 497830 258316 497836
rect 258172 456136 258224 456142
rect 258172 456078 258224 456084
rect 258080 452260 258132 452266
rect 258080 452202 258132 452208
rect 257448 449942 257738 449970
rect 258092 449956 258120 452202
rect 258276 449970 258304 497830
rect 258540 456136 258592 456142
rect 258540 456078 258592 456084
rect 258552 449970 258580 456078
rect 259184 452396 259236 452402
rect 259184 452338 259236 452344
rect 258276 449942 258474 449970
rect 258552 449942 258842 449970
rect 259196 449956 259224 452338
rect 259472 450158 259500 497898
rect 259460 450152 259512 450158
rect 259460 450094 259512 450100
rect 259564 449956 259592 497898
rect 259656 449970 259684 498034
rect 259734 495000 259790 495009
rect 259734 494935 259790 494944
rect 259748 460934 259776 494935
rect 259748 460906 260420 460934
rect 260012 450152 260064 450158
rect 260012 450094 260064 450100
rect 260024 449970 260052 450094
rect 260392 449970 260420 460906
rect 259656 449942 259946 449970
rect 260024 449942 260314 449970
rect 260392 449942 260682 449970
rect 261036 449956 261064 498918
rect 277398 496088 277454 496097
rect 277398 496023 277454 496032
rect 273352 464228 273404 464234
rect 273352 464170 273404 464176
rect 271880 464160 271932 464166
rect 271880 464102 271932 464108
rect 270776 464024 270828 464030
rect 270776 463966 270828 463972
rect 270592 461440 270644 461446
rect 270592 461382 270644 461388
rect 266360 461372 266412 461378
rect 266360 461314 266412 461320
rect 262956 458992 263008 458998
rect 262956 458934 263008 458940
rect 262588 454844 262640 454850
rect 262588 454786 262640 454792
rect 262128 453008 262180 453014
rect 262128 452950 262180 452956
rect 261760 452940 261812 452946
rect 261760 452882 261812 452888
rect 261772 449956 261800 452882
rect 262140 449956 262168 452950
rect 262220 452804 262272 452810
rect 262220 452746 262272 452752
rect 262232 449970 262260 452746
rect 262600 449970 262628 454786
rect 262968 449970 262996 458934
rect 264980 457292 265032 457298
rect 264980 457234 265032 457240
rect 264060 454776 264112 454782
rect 264060 454718 264112 454724
rect 263968 452736 264020 452742
rect 263968 452678 264020 452684
rect 262232 449942 262522 449970
rect 262600 449942 262890 449970
rect 262968 449942 263258 449970
rect 263980 449956 264008 452678
rect 264072 449970 264100 454718
rect 264702 452024 264758 452033
rect 264702 451959 264758 451968
rect 264072 449942 264362 449970
rect 264716 449956 264744 451959
rect 264992 449970 265020 457234
rect 265438 453248 265494 453257
rect 265438 453183 265494 453192
rect 264992 449942 265098 449970
rect 265452 449956 265480 453183
rect 265808 452872 265860 452878
rect 265808 452814 265860 452820
rect 265820 449956 265848 452814
rect 266174 451888 266230 451897
rect 266174 451823 266230 451832
rect 266188 449956 266216 451823
rect 266372 449970 266400 461314
rect 267740 461168 267792 461174
rect 267740 461110 267792 461116
rect 267004 458788 267056 458794
rect 267004 458730 267056 458736
rect 266910 451752 266966 451761
rect 266910 451687 266966 451696
rect 266372 449942 266570 449970
rect 266924 449956 266952 451687
rect 267016 449970 267044 458730
rect 267752 449970 267780 461110
rect 269120 459944 269172 459950
rect 269120 459886 269172 459892
rect 268108 454640 268160 454646
rect 268108 454582 268160 454588
rect 268120 449970 268148 454582
rect 267016 449942 267306 449970
rect 267752 449942 268042 449970
rect 268120 449942 268410 449970
rect 269132 449956 269160 459886
rect 269948 456340 270000 456346
rect 269948 456282 270000 456288
rect 269856 450492 269908 450498
rect 269856 450434 269908 450440
rect 269488 450424 269540 450430
rect 269488 450366 269540 450372
rect 269500 449956 269528 450366
rect 269868 449956 269896 450434
rect 269960 449970 269988 456282
rect 269960 449942 270250 449970
rect 270604 449956 270632 461382
rect 270684 461304 270736 461310
rect 270684 461246 270736 461252
rect 270696 456142 270724 461246
rect 270788 460934 270816 463966
rect 270788 460906 271092 460934
rect 270684 456136 270736 456142
rect 270684 456078 270736 456084
rect 270960 452668 271012 452674
rect 270960 452610 271012 452616
rect 270972 449956 271000 452610
rect 271064 449970 271092 460906
rect 271892 456142 271920 464102
rect 271972 464092 272024 464098
rect 271972 464034 272024 464040
rect 271420 456136 271472 456142
rect 271420 456078 271472 456084
rect 271880 456136 271932 456142
rect 271880 456078 271932 456084
rect 271432 449970 271460 456078
rect 271984 449970 272012 464034
rect 273258 463720 273314 463729
rect 273258 463655 273314 463664
rect 272154 461408 272210 461417
rect 272154 461343 272210 461352
rect 272064 461236 272116 461242
rect 272064 461178 272116 461184
rect 272076 451274 272104 461178
rect 272168 460934 272196 461343
rect 272168 460906 272932 460934
rect 272524 456136 272576 456142
rect 272524 456078 272576 456084
rect 272076 451246 272196 451274
rect 272168 449970 272196 451246
rect 272536 449970 272564 456078
rect 272904 449970 272932 460906
rect 273272 456142 273300 463655
rect 273260 456136 273312 456142
rect 273260 456078 273312 456084
rect 273364 449970 273392 464170
rect 274732 463956 274784 463962
rect 274732 463898 274784 463904
rect 273996 456136 274048 456142
rect 273996 456078 274048 456084
rect 273902 453112 273958 453121
rect 273902 453047 273958 453056
rect 271064 449942 271354 449970
rect 271432 449942 271722 449970
rect 271984 449942 272090 449970
rect 272168 449942 272458 449970
rect 272536 449942 272826 449970
rect 272904 449942 273194 449970
rect 273364 449942 273562 449970
rect 273916 449956 273944 453047
rect 274008 449970 274036 456078
rect 274744 449970 274772 463898
rect 274824 463888 274876 463894
rect 274824 463830 274876 463836
rect 274836 460934 274864 463830
rect 276204 463820 276256 463826
rect 276204 463762 276256 463768
rect 274836 460906 275140 460934
rect 275008 452124 275060 452130
rect 275008 452066 275060 452072
rect 274008 449942 274298 449970
rect 274666 449942 274772 449970
rect 275020 449956 275048 452066
rect 275112 449970 275140 460906
rect 276112 459876 276164 459882
rect 276112 459818 276164 459824
rect 275744 451784 275796 451790
rect 275744 451726 275796 451732
rect 275112 449942 275402 449970
rect 275756 449956 275784 451726
rect 276124 450430 276152 459818
rect 276112 450424 276164 450430
rect 276112 450366 276164 450372
rect 276216 449970 276244 463762
rect 277412 456142 277440 496023
rect 278044 495508 278096 495514
rect 278044 495450 278096 495456
rect 278056 465050 278084 495450
rect 286324 495236 286376 495242
rect 286324 495178 286376 495184
rect 280252 493536 280304 493542
rect 280252 493478 280304 493484
rect 280158 493368 280214 493377
rect 280158 493303 280214 493312
rect 278780 479664 278832 479670
rect 278780 479606 278832 479612
rect 277492 465044 277544 465050
rect 277492 464986 277544 464992
rect 278044 465044 278096 465050
rect 278044 464986 278096 464992
rect 277504 460934 277532 464986
rect 278792 460934 278820 479606
rect 277504 460906 278084 460934
rect 278792 460906 279188 460934
rect 277584 458720 277636 458726
rect 277584 458662 277636 458668
rect 277400 456136 277452 456142
rect 277400 456078 277452 456084
rect 277216 452192 277268 452198
rect 277216 452134 277268 452140
rect 276480 452056 276532 452062
rect 276480 451998 276532 452004
rect 276138 449942 276244 449970
rect 276492 449956 276520 451998
rect 276572 450424 276624 450430
rect 276572 450366 276624 450372
rect 276584 449970 276612 450366
rect 276584 449942 276874 449970
rect 277228 449956 277256 452134
rect 277596 449956 277624 458662
rect 277674 454744 277730 454753
rect 277674 454679 277730 454688
rect 277688 449970 277716 454679
rect 278056 449970 278084 460906
rect 278412 456136 278464 456142
rect 278412 456078 278464 456084
rect 278424 449970 278452 456078
rect 279056 452736 279108 452742
rect 279056 452678 279108 452684
rect 277688 449942 277978 449970
rect 278056 449942 278346 449970
rect 278424 449942 278714 449970
rect 279068 449956 279096 452678
rect 279160 449970 279188 460906
rect 279516 456272 279568 456278
rect 279516 456214 279568 456220
rect 279528 449970 279556 456214
rect 280172 456142 280200 493303
rect 280160 456136 280212 456142
rect 280160 456078 280212 456084
rect 280264 449970 280292 493478
rect 281816 490748 281868 490754
rect 281816 490690 281868 490696
rect 280804 489252 280856 489258
rect 280804 489194 280856 489200
rect 280620 456136 280672 456142
rect 280620 456078 280672 456084
rect 280528 453688 280580 453694
rect 280528 453630 280580 453636
rect 279160 449942 279450 449970
rect 279528 449942 279818 449970
rect 280186 449942 280292 449970
rect 280540 449956 280568 453630
rect 280632 449970 280660 456078
rect 280816 455938 280844 489194
rect 281828 484362 281856 490690
rect 286336 487150 286364 495178
rect 287060 489252 287112 489258
rect 287060 489194 287112 489200
rect 286324 487144 286376 487150
rect 286324 487086 286376 487092
rect 282920 486668 282972 486674
rect 282920 486610 282972 486616
rect 281816 484356 281868 484362
rect 281816 484298 281868 484304
rect 281724 465792 281776 465798
rect 281724 465734 281776 465740
rect 281632 463344 281684 463350
rect 281632 463286 281684 463292
rect 280988 459808 281040 459814
rect 280988 459750 281040 459756
rect 280804 455932 280856 455938
rect 280804 455874 280856 455880
rect 280816 452606 280844 455874
rect 280804 452600 280856 452606
rect 280804 452542 280856 452548
rect 281000 449970 281028 459750
rect 280632 449942 280922 449970
rect 281000 449942 281290 449970
rect 281644 449956 281672 463286
rect 281736 462398 281764 465734
rect 281724 462392 281776 462398
rect 281724 462334 281776 462340
rect 281736 456142 281764 462334
rect 281828 460934 281856 484298
rect 282932 460934 282960 486610
rect 286336 485926 286364 487086
rect 285680 485920 285732 485926
rect 285680 485862 285732 485868
rect 286324 485920 286376 485926
rect 286324 485862 286376 485868
rect 284484 468648 284536 468654
rect 284484 468590 284536 468596
rect 284496 460934 284524 468590
rect 281828 460906 282132 460934
rect 282932 460906 283604 460934
rect 284496 460906 285076 460934
rect 281724 456136 281776 456142
rect 281724 456078 281776 456084
rect 282000 452600 282052 452606
rect 282000 452542 282052 452548
rect 282012 449956 282040 452542
rect 282104 449970 282132 460906
rect 283010 456920 283066 456929
rect 283010 456855 283066 456864
rect 282460 456136 282512 456142
rect 282460 456078 282512 456084
rect 282472 449970 282500 456078
rect 283024 449970 283052 456855
rect 283472 452804 283524 452810
rect 283472 452746 283524 452752
rect 282104 449942 282394 449970
rect 282472 449942 282762 449970
rect 283024 449942 283130 449970
rect 283484 449956 283512 452746
rect 283576 449970 283604 460906
rect 284576 453552 284628 453558
rect 284576 453494 284628 453500
rect 284206 451616 284262 451625
rect 284206 451551 284262 451560
rect 283576 449942 283866 449970
rect 284220 449956 284248 451551
rect 284588 449956 284616 453494
rect 284942 453112 284998 453121
rect 284942 453047 284998 453056
rect 284956 449956 284984 453047
rect 285048 449970 285076 460906
rect 285692 456142 285720 485862
rect 285772 463276 285824 463282
rect 285772 463218 285824 463224
rect 285680 456136 285732 456142
rect 285680 456078 285732 456084
rect 285784 450430 285812 463218
rect 285864 463072 285916 463078
rect 285864 463014 285916 463020
rect 285876 456278 285904 463014
rect 285954 457600 286010 457609
rect 285954 457535 286010 457544
rect 285864 456272 285916 456278
rect 285864 456214 285916 456220
rect 285772 450424 285824 450430
rect 285772 450366 285824 450372
rect 285048 449942 285338 449970
rect 233422 449919 233478 449928
rect 225512 449890 225564 449896
rect 193864 449822 193916 449828
rect 219466 449806 219756 449834
rect 230478 449848 230534 449857
rect 285968 449834 285996 457535
rect 287072 456278 287100 489194
rect 287152 475516 287204 475522
rect 287152 475458 287204 475464
rect 287164 460934 287192 475458
rect 287702 474056 287758 474065
rect 287702 473991 287758 474000
rect 287716 465050 287744 473991
rect 287704 465044 287756 465050
rect 287704 464986 287756 464992
rect 288348 465044 288400 465050
rect 288348 464986 288400 464992
rect 287164 460906 287284 460934
rect 286140 456272 286192 456278
rect 286140 456214 286192 456220
rect 286600 456272 286652 456278
rect 286600 456214 286652 456220
rect 287060 456272 287112 456278
rect 287060 456214 287112 456220
rect 286048 450424 286100 450430
rect 286048 450366 286100 450372
rect 286060 449956 286088 450366
rect 286152 449970 286180 456214
rect 286612 456142 286640 456214
rect 286508 456136 286560 456142
rect 286508 456078 286560 456084
rect 286600 456136 286652 456142
rect 286600 456078 286652 456084
rect 286520 449970 286548 456078
rect 287152 452532 287204 452538
rect 287152 452474 287204 452480
rect 286152 449942 286442 449970
rect 286520 449942 286810 449970
rect 287164 449956 287192 452474
rect 287256 449970 287284 460906
rect 287980 456272 288032 456278
rect 287980 456214 288032 456220
rect 287886 451344 287942 451353
rect 287886 451279 287942 451288
rect 287256 449942 287546 449970
rect 287900 449956 287928 451279
rect 287992 449970 288020 456214
rect 288360 452538 288388 464986
rect 288452 456278 288480 500375
rect 302240 498160 302292 498166
rect 302240 498102 302292 498108
rect 301504 496936 301556 496942
rect 301504 496878 301556 496884
rect 293960 493468 294012 493474
rect 293960 493410 294012 493416
rect 293972 492726 294000 493410
rect 293960 492720 294012 492726
rect 293960 492662 294012 492668
rect 294236 492720 294288 492726
rect 294236 492662 294288 492668
rect 292488 490884 292540 490890
rect 292488 490826 292540 490832
rect 291200 489864 291252 489870
rect 291200 489806 291252 489812
rect 291212 488782 291240 489806
rect 292500 488782 292528 490826
rect 291200 488776 291252 488782
rect 291200 488718 291252 488724
rect 292488 488776 292540 488782
rect 292488 488718 292540 488724
rect 290464 474156 290516 474162
rect 290464 474098 290516 474104
rect 288532 471300 288584 471306
rect 288532 471242 288584 471248
rect 288544 460934 288572 471242
rect 290476 464506 290504 474098
rect 290464 464500 290516 464506
rect 290464 464442 290516 464448
rect 290476 464234 290504 464442
rect 289820 464228 289872 464234
rect 289820 464170 289872 464176
rect 290464 464228 290516 464234
rect 290464 464170 290516 464176
rect 289832 460934 289860 464170
rect 288544 460906 288756 460934
rect 289832 460906 290596 460934
rect 288440 456272 288492 456278
rect 288440 456214 288492 456220
rect 288348 452532 288400 452538
rect 288348 452474 288400 452480
rect 288624 450356 288676 450362
rect 288624 450298 288676 450304
rect 287992 449942 288282 449970
rect 288636 449956 288664 450298
rect 288728 449970 288756 460906
rect 290188 460624 290240 460630
rect 290188 460566 290240 460572
rect 289452 456272 289504 456278
rect 289452 456214 289504 456220
rect 290002 456240 290058 456249
rect 289082 454336 289138 454345
rect 289082 454271 289138 454280
rect 289096 449970 289124 454271
rect 289464 449970 289492 456214
rect 290002 456175 290058 456184
rect 290016 449970 290044 456175
rect 290200 449970 290228 460566
rect 290568 449970 290596 460906
rect 288728 449942 289018 449970
rect 289096 449942 289386 449970
rect 289464 449942 289754 449970
rect 290016 449942 290122 449970
rect 290200 449942 290490 449970
rect 290568 449942 290858 449970
rect 291212 449956 291240 488718
rect 292856 488028 292908 488034
rect 292856 487970 292908 487976
rect 291292 467152 291344 467158
rect 291292 467094 291344 467100
rect 291304 465186 291332 467094
rect 291292 465180 291344 465186
rect 291292 465122 291344 465128
rect 291304 449970 291332 465122
rect 291936 452940 291988 452946
rect 291936 452882 291988 452888
rect 291304 449942 291594 449970
rect 291948 449956 291976 452882
rect 292302 451616 292358 451625
rect 292302 451551 292358 451560
rect 292316 449956 292344 451551
rect 292868 449970 292896 487970
rect 294052 474156 294104 474162
rect 294052 474098 294104 474104
rect 293040 456408 293092 456414
rect 293040 456350 293092 456356
rect 292698 449942 292896 449970
rect 293052 449956 293080 456350
rect 293776 454164 293828 454170
rect 293776 454106 293828 454112
rect 293408 453484 293460 453490
rect 293408 453426 293460 453432
rect 293420 449956 293448 453426
rect 293788 449956 293816 454106
rect 294064 449970 294092 474098
rect 294248 466454 294276 492662
rect 301044 490748 301096 490754
rect 301044 490690 301096 490696
rect 300124 487892 300176 487898
rect 300124 487834 300176 487840
rect 296904 483812 296956 483818
rect 296904 483754 296956 483760
rect 295340 478236 295392 478242
rect 295340 478178 295392 478184
rect 294248 466426 295012 466454
rect 294144 461100 294196 461106
rect 294144 461042 294196 461048
rect 294156 456794 294184 461042
rect 294604 460556 294656 460562
rect 294604 460498 294656 460504
rect 294156 456766 294276 456794
rect 294248 449970 294276 456766
rect 294616 449970 294644 460498
rect 294984 449970 295012 466426
rect 295352 453014 295380 478178
rect 295432 468512 295484 468518
rect 295432 468454 295484 468460
rect 295444 466546 295472 468454
rect 295432 466540 295484 466546
rect 295432 466482 295484 466488
rect 295444 453082 295472 466482
rect 295708 465112 295760 465118
rect 295708 465054 295760 465060
rect 295720 462466 295748 465054
rect 295708 462460 295760 462466
rect 295708 462402 295760 462408
rect 295432 453076 295484 453082
rect 295432 453018 295484 453024
rect 295340 453008 295392 453014
rect 295340 452950 295392 452956
rect 295720 449970 295748 462402
rect 295800 453076 295852 453082
rect 295800 453018 295852 453024
rect 294064 449942 294170 449970
rect 294248 449942 294538 449970
rect 294616 449942 294906 449970
rect 294984 449942 295274 449970
rect 295642 449942 295748 449970
rect 295812 449970 295840 453018
rect 296076 453008 296128 453014
rect 296076 452950 296128 452956
rect 296088 449970 296116 452950
rect 296720 451716 296772 451722
rect 296720 451658 296772 451664
rect 295812 449942 296010 449970
rect 296088 449942 296378 449970
rect 296732 449956 296760 451658
rect 296916 449970 296944 483754
rect 300136 468722 300164 487834
rect 300768 469872 300820 469878
rect 300768 469814 300820 469820
rect 300780 469198 300808 469814
rect 300768 469192 300820 469198
rect 300768 469134 300820 469140
rect 300124 468716 300176 468722
rect 300124 468658 300176 468664
rect 300136 467906 300164 468658
rect 299480 467900 299532 467906
rect 299480 467842 299532 467848
rect 300124 467900 300176 467906
rect 300124 467842 300176 467848
rect 298284 461712 298336 461718
rect 298284 461654 298336 461660
rect 297824 453416 297876 453422
rect 297824 453358 297876 453364
rect 297456 450220 297508 450226
rect 297456 450162 297508 450168
rect 296916 449942 297114 449970
rect 297468 449956 297496 450162
rect 297836 449956 297864 453358
rect 298192 452872 298244 452878
rect 298192 452814 298244 452820
rect 298204 449956 298232 452814
rect 298296 449970 298324 461654
rect 299020 460488 299072 460494
rect 299020 460430 299072 460436
rect 298926 450664 298982 450673
rect 298926 450599 298982 450608
rect 298296 449942 298586 449970
rect 298940 449956 298968 450599
rect 299032 449970 299060 460430
rect 299492 449970 299520 467842
rect 300398 452840 300454 452849
rect 300398 452775 300454 452784
rect 300032 452396 300084 452402
rect 300032 452338 300084 452344
rect 299032 449942 299322 449970
rect 299492 449942 299690 449970
rect 300044 449956 300072 452338
rect 300412 449956 300440 452775
rect 300780 452402 300808 469134
rect 300768 452396 300820 452402
rect 300768 452338 300820 452344
rect 300766 451888 300822 451897
rect 300766 451823 300822 451832
rect 300780 449956 300808 451823
rect 301056 449970 301084 490690
rect 301516 480282 301544 496878
rect 301504 480276 301556 480282
rect 301504 480218 301556 480224
rect 301516 465798 301544 480218
rect 301504 465792 301556 465798
rect 301504 465734 301556 465740
rect 301228 459740 301280 459746
rect 301228 459682 301280 459688
rect 301240 449970 301268 459682
rect 301872 453348 301924 453354
rect 301872 453290 301924 453296
rect 301056 449942 301162 449970
rect 301240 449942 301530 449970
rect 301884 449956 301912 453290
rect 302252 450362 302280 498102
rect 313280 497480 313332 497486
rect 313280 497422 313332 497428
rect 313292 497010 313320 497422
rect 319444 497072 319496 497078
rect 319444 497014 319496 497020
rect 313280 497004 313332 497010
rect 313280 496946 313332 496952
rect 315304 497004 315356 497010
rect 315304 496946 315356 496952
rect 311164 496936 311216 496942
rect 311164 496878 311216 496884
rect 305000 496120 305052 496126
rect 305000 496062 305052 496068
rect 304356 494828 304408 494834
rect 304356 494770 304408 494776
rect 303804 474224 303856 474230
rect 303804 474166 303856 474172
rect 303712 469260 303764 469266
rect 303712 469202 303764 469208
rect 302330 463040 302386 463049
rect 302330 462975 302386 462984
rect 302344 460934 302372 462975
rect 302344 460906 302740 460934
rect 302516 458720 302568 458726
rect 302516 458662 302568 458668
rect 302240 450356 302292 450362
rect 302240 450298 302292 450304
rect 302528 449834 302556 458662
rect 302608 450356 302660 450362
rect 302608 450298 302660 450304
rect 302620 449956 302648 450298
rect 302712 449970 302740 460906
rect 303068 460420 303120 460426
rect 303068 460362 303120 460368
rect 303080 449970 303108 460362
rect 303620 456272 303672 456278
rect 303620 456214 303672 456220
rect 303632 449970 303660 456214
rect 303724 451274 303752 469202
rect 303816 460934 303844 474166
rect 304368 469266 304396 494770
rect 304356 469260 304408 469266
rect 304356 469202 304408 469208
rect 304264 465792 304316 465798
rect 304264 465734 304316 465740
rect 303816 460906 304212 460934
rect 303724 451246 303844 451274
rect 303816 449970 303844 451246
rect 304184 449970 304212 460906
rect 304276 456278 304304 465734
rect 305012 456278 305040 496062
rect 305092 482520 305144 482526
rect 305092 482462 305144 482468
rect 304264 456272 304316 456278
rect 304264 456214 304316 456220
rect 305000 456272 305052 456278
rect 305000 456214 305052 456220
rect 304814 449984 304870 449993
rect 302712 449942 303002 449970
rect 303080 449942 303370 449970
rect 303632 449942 303738 449970
rect 303816 449942 304106 449970
rect 304184 449942 304474 449970
rect 305104 449970 305132 482462
rect 309140 481092 309192 481098
rect 309140 481034 309192 481040
rect 307024 476944 307076 476950
rect 307024 476886 307076 476892
rect 307036 469402 307064 476886
rect 308496 472660 308548 472666
rect 308496 472602 308548 472608
rect 307024 469396 307076 469402
rect 307024 469338 307076 469344
rect 306380 461032 306432 461038
rect 306380 460974 306432 460980
rect 306392 460934 306420 460974
rect 306392 460906 306788 460934
rect 306012 458788 306064 458794
rect 306012 458730 306064 458736
rect 305644 456272 305696 456278
rect 305644 456214 305696 456220
rect 305552 450288 305604 450294
rect 305552 450230 305604 450236
rect 305104 449942 305210 449970
rect 305564 449956 305592 450230
rect 305656 449970 305684 456214
rect 306024 449970 306052 458730
rect 306656 452056 306708 452062
rect 306656 451998 306708 452004
rect 305656 449942 305946 449970
rect 306024 449942 306314 449970
rect 306668 449956 306696 451998
rect 306760 449970 306788 460906
rect 307036 452606 307064 469338
rect 308508 463690 308536 472602
rect 308496 463684 308548 463690
rect 308496 463626 308548 463632
rect 309048 463684 309100 463690
rect 309048 463626 309100 463632
rect 307116 460352 307168 460358
rect 307116 460294 307168 460300
rect 307024 452600 307076 452606
rect 307024 452542 307076 452548
rect 307128 449970 307156 460294
rect 309060 452606 309088 463626
rect 308036 452600 308088 452606
rect 308036 452542 308088 452548
rect 308128 452600 308180 452606
rect 308128 452542 308180 452548
rect 309048 452600 309100 452606
rect 309048 452542 309100 452548
rect 308048 449970 308076 452542
rect 308140 451382 308168 452542
rect 308496 452328 308548 452334
rect 308496 452270 308548 452276
rect 308128 451376 308180 451382
rect 308128 451318 308180 451324
rect 306760 449942 307050 449970
rect 307128 449942 307418 449970
rect 307786 449942 308076 449970
rect 308140 449956 308168 451318
rect 308508 449956 308536 452270
rect 309152 449970 309180 481034
rect 309232 481024 309284 481030
rect 309232 480966 309284 480972
rect 309244 460934 309272 480966
rect 311176 470558 311204 496878
rect 313280 490680 313332 490686
rect 313280 490622 313332 490628
rect 311900 476808 311952 476814
rect 311900 476750 311952 476756
rect 311912 472054 311940 476750
rect 311900 472048 311952 472054
rect 311900 471990 311952 471996
rect 311164 470552 311216 470558
rect 311164 470494 311216 470500
rect 311176 469334 311204 470494
rect 310520 469328 310572 469334
rect 310520 469270 310572 469276
rect 311164 469328 311216 469334
rect 311164 469270 311216 469276
rect 309244 460906 309732 460934
rect 309322 458960 309378 458969
rect 309322 458895 309378 458904
rect 309336 449970 309364 458895
rect 309704 449970 309732 460906
rect 310060 458652 310112 458658
rect 310060 458594 310112 458600
rect 310072 449970 310100 458594
rect 310532 456346 310560 469270
rect 310612 465860 310664 465866
rect 310612 465802 310664 465808
rect 310520 456340 310572 456346
rect 310520 456282 310572 456288
rect 310624 456278 310652 465802
rect 310702 462768 310758 462777
rect 310702 462703 310758 462712
rect 310716 460934 310744 462703
rect 310716 460906 310836 460934
rect 310612 456272 310664 456278
rect 310612 456214 310664 456220
rect 310704 452124 310756 452130
rect 310704 452066 310756 452072
rect 309152 449942 309258 449970
rect 309336 449942 309626 449970
rect 309704 449942 309994 449970
rect 310072 449942 310362 449970
rect 310716 449956 310744 452066
rect 310808 449970 310836 460906
rect 311532 456340 311584 456346
rect 311532 456282 311584 456288
rect 311164 456272 311216 456278
rect 311164 456214 311216 456220
rect 311176 449970 311204 456214
rect 311544 449970 311572 456282
rect 311912 449970 311940 471990
rect 311992 471300 312044 471306
rect 311992 471242 312044 471248
rect 312004 460934 312032 471242
rect 312004 460906 312676 460934
rect 312648 449970 312676 460906
rect 313188 458516 313240 458522
rect 313188 458458 313240 458464
rect 313200 458130 313228 458458
rect 313292 458266 313320 490622
rect 313372 467288 313424 467294
rect 313372 467230 313424 467236
rect 313384 460934 313412 467230
rect 314658 466032 314714 466041
rect 314658 465967 314714 465976
rect 313384 460906 314148 460934
rect 313740 458584 313792 458590
rect 313740 458526 313792 458532
rect 313292 458238 313412 458266
rect 313200 458102 313320 458130
rect 310808 449942 311098 449970
rect 311176 449942 311466 449970
rect 311544 449942 311834 449970
rect 311912 449942 312202 449970
rect 312648 449942 312938 449970
rect 313292 449956 313320 458102
rect 313384 449970 313412 458238
rect 313752 449970 313780 458526
rect 314120 449970 314148 460906
rect 313384 449942 313674 449970
rect 313752 449942 314042 449970
rect 314120 449942 314410 449970
rect 314672 449954 314700 465967
rect 314750 461272 314806 461281
rect 314750 461207 314806 461216
rect 314764 460934 314792 461207
rect 314764 460906 314976 460934
rect 314948 450106 314976 460906
rect 315316 451274 315344 496946
rect 316040 496120 316092 496126
rect 316040 496062 316092 496068
rect 315856 453076 315908 453082
rect 315856 453018 315908 453024
rect 314764 450078 314976 450106
rect 315224 451246 315344 451274
rect 314764 449956 314792 450078
rect 315224 449970 315252 451246
rect 314948 449954 315146 449970
rect 314660 449948 314712 449954
rect 304814 449919 304870 449928
rect 314660 449890 314712 449896
rect 314936 449948 315146 449954
rect 314988 449942 315146 449948
rect 315224 449942 315514 449970
rect 315868 449956 315896 453018
rect 316052 449970 316080 496062
rect 319076 494828 319128 494834
rect 319076 494770 319128 494776
rect 316132 482452 316184 482458
rect 316132 482394 316184 482400
rect 316144 460934 316172 482394
rect 318892 478916 318944 478922
rect 318892 478858 318944 478864
rect 317418 465896 317474 465905
rect 317418 465831 317474 465840
rect 316144 460906 316724 460934
rect 316590 450528 316646 450537
rect 316590 450463 316646 450472
rect 316052 449942 316250 449970
rect 316604 449956 316632 450463
rect 316696 449970 316724 460906
rect 317052 458516 317104 458522
rect 317052 458458 317104 458464
rect 317064 449970 317092 458458
rect 317328 456272 317380 456278
rect 317328 456214 317380 456220
rect 317340 456006 317368 456214
rect 317432 456006 317460 465831
rect 317510 462632 317566 462641
rect 317510 462567 317566 462576
rect 317524 460934 317552 462567
rect 317524 460906 317828 460934
rect 317328 456000 317380 456006
rect 317328 455942 317380 455948
rect 317420 456000 317472 456006
rect 317420 455942 317472 455948
rect 317696 452192 317748 452198
rect 317696 452134 317748 452140
rect 316696 449942 316986 449970
rect 317064 449942 317354 449970
rect 317708 449956 317736 452134
rect 317800 449970 317828 460906
rect 318156 456000 318208 456006
rect 318156 455942 318208 455948
rect 318168 449970 318196 455942
rect 318904 449970 318932 478858
rect 319088 460934 319116 494770
rect 319456 480214 319484 497014
rect 319444 480208 319496 480214
rect 319444 480150 319496 480156
rect 319456 478922 319484 480150
rect 319444 478916 319496 478922
rect 319444 478858 319496 478864
rect 319088 460906 319300 460934
rect 319166 451752 319222 451761
rect 319166 451687 319222 451696
rect 317800 449942 318090 449970
rect 318168 449942 318458 449970
rect 318826 449942 318932 449970
rect 319180 449956 319208 451687
rect 319272 449970 319300 460906
rect 319628 457224 319680 457230
rect 319628 457166 319680 457172
rect 319640 449970 319668 457166
rect 320192 456006 320220 500511
rect 336740 500482 336792 500488
rect 333980 500472 334032 500478
rect 333980 500414 334032 500420
rect 329840 500404 329892 500410
rect 329840 500346 329892 500352
rect 327080 500336 327132 500342
rect 327080 500278 327132 500284
rect 324596 500268 324648 500274
rect 324596 500210 324648 500216
rect 320272 492040 320324 492046
rect 320272 491982 320324 491988
rect 320180 456000 320232 456006
rect 320180 455942 320232 455948
rect 319272 449942 319562 449970
rect 319640 449942 319930 449970
rect 320284 449956 320312 491982
rect 322940 490612 322992 490618
rect 322940 490554 322992 490560
rect 321560 476808 321612 476814
rect 321560 476750 321612 476756
rect 321100 459264 321152 459270
rect 321100 459206 321152 459212
rect 320732 456000 320784 456006
rect 320732 455942 320784 455948
rect 320638 450528 320694 450537
rect 320638 450463 320694 450472
rect 320652 449956 320680 450463
rect 320744 449970 320772 455942
rect 321112 449970 321140 459206
rect 321572 453014 321600 476750
rect 322204 475448 322256 475454
rect 322204 475390 322256 475396
rect 321652 467220 321704 467226
rect 321652 467162 321704 467168
rect 321560 453008 321612 453014
rect 321560 452950 321612 452956
rect 321664 449970 321692 467162
rect 322216 456346 322244 475390
rect 322952 456794 322980 490554
rect 324504 487212 324556 487218
rect 324504 487154 324556 487160
rect 324516 485790 324544 487154
rect 324504 485784 324556 485790
rect 324504 485726 324556 485732
rect 324516 480254 324544 485726
rect 324424 480226 324544 480254
rect 324320 459672 324372 459678
rect 324320 459614 324372 459620
rect 322952 456766 323348 456794
rect 322204 456340 322256 456346
rect 322204 456282 322256 456288
rect 322216 449970 322244 456282
rect 323216 456272 323268 456278
rect 323216 456214 323268 456220
rect 322572 453008 322624 453014
rect 322572 452950 322624 452956
rect 322480 451784 322532 451790
rect 322480 451726 322532 451732
rect 320744 449942 321034 449970
rect 321112 449942 321402 449970
rect 321664 449942 321770 449970
rect 322138 449942 322244 449970
rect 322492 449956 322520 451726
rect 322584 449970 322612 452950
rect 322584 449942 322874 449970
rect 323228 449956 323256 456214
rect 323320 449970 323348 456766
rect 323952 454232 324004 454238
rect 323952 454174 324004 454180
rect 323320 449942 323610 449970
rect 323964 449956 323992 454174
rect 324332 453218 324360 459614
rect 324320 453212 324372 453218
rect 324320 453154 324372 453160
rect 324424 453014 324452 480226
rect 324504 472864 324556 472870
rect 324504 472806 324556 472812
rect 324516 453150 324544 472806
rect 324504 453144 324556 453150
rect 324504 453086 324556 453092
rect 324412 453008 324464 453014
rect 324412 452950 324464 452956
rect 314936 449890 314988 449896
rect 324608 449834 324636 500210
rect 325976 493468 326028 493474
rect 325976 493410 326028 493416
rect 325792 489184 325844 489190
rect 325792 489126 325844 489132
rect 324688 453212 324740 453218
rect 324688 453154 324740 453160
rect 324700 449956 324728 453154
rect 324780 453144 324832 453150
rect 324780 453086 324832 453092
rect 324792 449970 324820 453086
rect 325804 453014 325832 489126
rect 325148 453008 325200 453014
rect 325148 452950 325200 452956
rect 325792 453008 325844 453014
rect 325792 452950 325844 452956
rect 325160 449970 325188 452950
rect 325792 452668 325844 452674
rect 325792 452610 325844 452616
rect 324792 449942 325082 449970
rect 325160 449942 325450 449970
rect 325804 449956 325832 452610
rect 325988 449970 326016 493410
rect 326252 457156 326304 457162
rect 326252 457098 326304 457104
rect 326264 449970 326292 457098
rect 327092 456794 327120 500278
rect 328460 492040 328512 492046
rect 328460 491982 328512 491988
rect 327172 483880 327224 483886
rect 327172 483822 327224 483828
rect 327184 460934 327212 483822
rect 327184 460906 328132 460934
rect 327724 459196 327776 459202
rect 327724 459138 327776 459144
rect 327092 456766 327396 456794
rect 327264 454300 327316 454306
rect 327264 454242 327316 454248
rect 326620 453008 326672 453014
rect 326620 452950 326672 452956
rect 326632 449970 326660 452950
rect 325988 449942 326186 449970
rect 326264 449942 326554 449970
rect 326632 449942 326922 449970
rect 327276 449956 327304 454242
rect 327368 449970 327396 456766
rect 327736 449970 327764 459138
rect 328104 449970 328132 460906
rect 328472 453014 328500 491982
rect 329104 491360 329156 491366
rect 329104 491302 329156 491308
rect 329116 471986 329144 491302
rect 328552 471980 328604 471986
rect 328552 471922 328604 471928
rect 329104 471980 329156 471986
rect 329104 471922 329156 471928
rect 328460 453008 328512 453014
rect 328460 452950 328512 452956
rect 328564 449970 328592 471922
rect 329852 453014 329880 500346
rect 332600 482384 332652 482390
rect 332600 482326 332652 482332
rect 329932 480956 329984 480962
rect 329932 480898 329984 480904
rect 329196 453008 329248 453014
rect 329196 452950 329248 452956
rect 329840 453008 329892 453014
rect 329840 452950 329892 452956
rect 329104 450220 329156 450226
rect 329104 450162 329156 450168
rect 327368 449942 327658 449970
rect 327736 449942 328026 449970
rect 328104 449942 328394 449970
rect 328564 449942 328762 449970
rect 329116 449956 329144 450162
rect 329208 449970 329236 452950
rect 329838 450392 329894 450401
rect 329838 450327 329894 450336
rect 329208 449942 329498 449970
rect 329852 449956 329880 450327
rect 329944 449970 329972 480898
rect 331220 472728 331272 472734
rect 331220 472670 331272 472676
rect 331232 471442 331260 472670
rect 331220 471436 331272 471442
rect 331220 471378 331272 471384
rect 331232 456006 331260 471378
rect 331312 468580 331364 468586
rect 331312 468522 331364 468528
rect 331324 460934 331352 468522
rect 331324 460906 331536 460934
rect 331402 460320 331458 460329
rect 331402 460255 331458 460264
rect 331220 456000 331272 456006
rect 331220 455942 331272 455948
rect 330576 453144 330628 453150
rect 330576 453086 330628 453092
rect 329944 449942 330234 449970
rect 330588 449956 330616 453086
rect 330668 453008 330720 453014
rect 330668 452950 330720 452956
rect 330760 453008 330812 453014
rect 330760 452950 330812 452956
rect 330680 449970 330708 452950
rect 330772 452674 330800 452950
rect 330760 452668 330812 452674
rect 330760 452610 330812 452616
rect 331416 449970 331444 460255
rect 330680 449942 330970 449970
rect 331338 449942 331444 449970
rect 331508 449970 331536 460906
rect 332612 456006 332640 482326
rect 332692 478236 332744 478242
rect 332692 478178 332744 478184
rect 331772 456000 331824 456006
rect 331772 455942 331824 455948
rect 332600 456000 332652 456006
rect 332600 455942 332652 455948
rect 331784 449970 331812 455942
rect 332416 450152 332468 450158
rect 332416 450094 332468 450100
rect 331508 449942 331706 449970
rect 331784 449942 332074 449970
rect 332428 449956 332456 450094
rect 332704 449970 332732 478178
rect 332874 456104 332930 456113
rect 332874 456039 332930 456048
rect 332888 449970 332916 456039
rect 333244 456000 333296 456006
rect 333244 455942 333296 455948
rect 333256 449970 333284 455942
rect 333612 454640 333664 454646
rect 333612 454582 333664 454588
rect 333624 449970 333652 454582
rect 333992 449970 334020 500414
rect 334912 497486 334940 500140
rect 334900 497480 334952 497486
rect 334900 497422 334952 497428
rect 334072 487960 334124 487966
rect 334072 487902 334124 487908
rect 334084 460934 334112 487902
rect 335360 480956 335412 480962
rect 335360 480898 335412 480904
rect 334084 460906 334756 460934
rect 334348 458448 334400 458454
rect 334348 458390 334400 458396
rect 334360 449970 334388 458390
rect 334728 449970 334756 460906
rect 335372 456006 335400 480898
rect 336648 465112 336700 465118
rect 336648 465054 336700 465060
rect 336660 463758 336688 465054
rect 335452 463752 335504 463758
rect 335452 463694 335504 463700
rect 336648 463752 336700 463758
rect 336648 463694 336700 463700
rect 335360 456000 335412 456006
rect 335360 455942 335412 455948
rect 335464 449970 335492 463694
rect 336752 456006 336780 500482
rect 340880 500200 340932 500206
rect 340880 500142 340932 500148
rect 338764 495576 338816 495582
rect 338764 495518 338816 495524
rect 336832 483744 336884 483750
rect 336832 483686 336884 483692
rect 335820 456000 335872 456006
rect 335820 455942 335872 455948
rect 336740 456000 336792 456006
rect 336740 455942 336792 455948
rect 335636 450084 335688 450090
rect 335636 450026 335688 450032
rect 332704 449942 332810 449970
rect 332888 449942 333178 449970
rect 333256 449942 333546 449970
rect 333624 449942 333914 449970
rect 333992 449942 334282 449970
rect 334360 449942 334650 449970
rect 334728 449942 335018 449970
rect 335386 449942 335492 449970
rect 335648 449970 335676 450026
rect 335832 449970 335860 455942
rect 336280 450016 336332 450022
rect 335648 449942 335754 449970
rect 335832 449942 336122 449970
rect 336332 449964 336490 449970
rect 336280 449958 336490 449964
rect 336292 449942 336490 449958
rect 336844 449956 336872 483686
rect 338120 482384 338172 482390
rect 338120 482326 338172 482332
rect 337658 460048 337714 460057
rect 337658 459983 337714 459992
rect 337292 456000 337344 456006
rect 337292 455942 337344 455948
rect 337200 453280 337252 453286
rect 337200 453222 337252 453228
rect 337212 449956 337240 453222
rect 337304 449970 337332 455942
rect 337672 449970 337700 459983
rect 338132 456006 338160 482326
rect 338210 475416 338266 475425
rect 338210 475351 338266 475360
rect 338120 456000 338172 456006
rect 338120 455942 338172 455948
rect 338224 449970 338252 475351
rect 338776 466478 338804 495518
rect 339500 487824 339552 487830
rect 339500 487766 339552 487772
rect 338304 466472 338356 466478
rect 338304 466414 338356 466420
rect 338764 466472 338816 466478
rect 338764 466414 338816 466420
rect 338316 460934 338344 466414
rect 339512 460934 339540 487766
rect 338316 460906 338436 460934
rect 339512 460906 339908 460934
rect 338408 449970 338436 460906
rect 339132 456000 339184 456006
rect 339132 455942 339184 455948
rect 338948 450016 339000 450022
rect 337304 449942 337594 449970
rect 337672 449942 337962 449970
rect 338224 449942 338330 449970
rect 338408 449942 338698 449970
rect 339144 449970 339172 455942
rect 339776 450900 339828 450906
rect 339776 450842 339828 450848
rect 339000 449964 339066 449970
rect 338948 449958 339066 449964
rect 338960 449942 339066 449958
rect 339144 449942 339434 449970
rect 339788 449956 339816 450842
rect 339880 449970 339908 460906
rect 340510 450392 340566 450401
rect 340510 450327 340566 450336
rect 339880 449942 340170 449970
rect 340524 449956 340552 450327
rect 340892 449956 340920 500142
rect 342260 490612 342312 490618
rect 342260 490554 342312 490560
rect 340972 479596 341024 479602
rect 340972 479538 341024 479544
rect 340984 460934 341012 479538
rect 340984 460906 341380 460934
rect 341064 458380 341116 458386
rect 341064 458322 341116 458328
rect 341076 449970 341104 458322
rect 341352 449970 341380 460906
rect 341984 450900 342036 450906
rect 341984 450842 342036 450848
rect 341076 449942 341274 449970
rect 341352 449942 341642 449970
rect 341996 449956 342024 450842
rect 342272 449970 342300 490554
rect 342352 486532 342404 486538
rect 342352 486474 342404 486480
rect 342364 460934 342392 486474
rect 342364 460906 342852 460934
rect 342534 457328 342590 457337
rect 342534 457263 342590 457272
rect 342548 449970 342576 457263
rect 342824 449970 342852 460906
rect 343180 454776 343232 454782
rect 343180 454718 343232 454724
rect 343192 449970 343220 454718
rect 343652 449970 343680 500550
rect 345020 483744 345072 483750
rect 345020 483686 345072 483692
rect 343732 471368 343784 471374
rect 343732 471310 343784 471316
rect 343744 460934 343772 471310
rect 343744 460906 344324 460934
rect 343914 459912 343970 459921
rect 343914 459847 343970 459856
rect 343928 449970 343956 459847
rect 344296 449970 344324 460906
rect 344928 453212 344980 453218
rect 344928 453154 344980 453160
rect 342272 449942 342378 449970
rect 342548 449942 342746 449970
rect 342824 449942 343114 449970
rect 343192 449942 343482 449970
rect 343652 449942 343850 449970
rect 343928 449942 344218 449970
rect 344296 449942 344586 449970
rect 344940 449956 344968 453154
rect 345032 449970 345060 483686
rect 345112 479528 345164 479534
rect 345112 479470 345164 479476
rect 345124 460934 345152 479470
rect 345124 460906 345796 460934
rect 345664 450968 345716 450974
rect 345664 450910 345716 450916
rect 345032 449942 345322 449970
rect 345676 449956 345704 450910
rect 345768 449970 345796 460906
rect 346412 458130 346440 500618
rect 349356 489914 349384 500686
rect 349620 500608 349672 500614
rect 349620 500550 349672 500556
rect 349632 500206 349660 500550
rect 351840 500206 351868 500686
rect 354956 500686 355008 500692
rect 364064 500744 364116 500750
rect 364156 500744 364208 500750
rect 364064 500686 364116 500692
rect 364154 500712 364156 500721
rect 364616 500744 364668 500750
rect 364208 500712 364210 500721
rect 354862 500647 354918 500656
rect 349620 500200 349672 500206
rect 349620 500142 349672 500148
rect 351828 500200 351880 500206
rect 351828 500142 351880 500148
rect 351920 500132 351972 500138
rect 351920 500074 351972 500080
rect 349172 489886 349384 489914
rect 346492 486600 346544 486606
rect 346492 486542 346544 486548
rect 346504 460934 346532 486542
rect 347780 485104 347832 485110
rect 347780 485046 347832 485052
rect 346504 460906 347268 460934
rect 346858 458824 346914 458833
rect 346858 458759 346914 458768
rect 346412 458102 346532 458130
rect 346400 453348 346452 453354
rect 346400 453290 346452 453296
rect 345768 449942 346058 449970
rect 346412 449956 346440 453290
rect 346504 449970 346532 458102
rect 346872 449970 346900 458759
rect 347240 449970 347268 460906
rect 347792 456006 347820 485046
rect 347872 461644 347924 461650
rect 347872 461586 347924 461592
rect 347884 460934 347912 461586
rect 347884 460906 348004 460934
rect 347780 456000 347832 456006
rect 347780 455942 347832 455948
rect 347872 450288 347924 450294
rect 347872 450230 347924 450236
rect 346504 449942 346794 449970
rect 346872 449942 347162 449970
rect 347240 449942 347530 449970
rect 347884 449956 347912 450230
rect 347976 449970 348004 460906
rect 348700 456000 348752 456006
rect 348330 455968 348386 455977
rect 348700 455942 348752 455948
rect 348330 455903 348386 455912
rect 348344 449970 348372 455903
rect 348712 449970 348740 455942
rect 349172 451274 349200 489886
rect 349252 489320 349304 489326
rect 349252 489262 349304 489268
rect 349264 460934 349292 489262
rect 350540 487824 350592 487830
rect 350540 487766 350592 487772
rect 350552 460934 350580 487766
rect 349264 460906 350212 460934
rect 350552 460906 350948 460934
rect 350078 452976 350134 452985
rect 350078 452911 350134 452920
rect 349172 451246 349476 451274
rect 349448 449970 349476 451246
rect 347976 449942 348266 449970
rect 348344 449942 348634 449970
rect 348712 449942 349002 449970
rect 349448 449942 349738 449970
rect 350092 449956 350120 452911
rect 350184 449970 350212 460906
rect 350816 450356 350868 450362
rect 350816 450298 350868 450304
rect 350184 449942 350474 449970
rect 350828 449956 350856 450298
rect 350920 449970 350948 460906
rect 351932 456006 351960 500074
rect 354968 495434 354996 500686
rect 357348 500200 357400 500206
rect 357348 500142 357400 500148
rect 357440 500200 357492 500206
rect 357440 500142 357492 500148
rect 357360 500070 357388 500142
rect 357348 500064 357400 500070
rect 357348 500006 357400 500012
rect 354692 495406 354996 495434
rect 353300 489184 353352 489190
rect 353300 489126 353352 489132
rect 352012 475380 352064 475386
rect 352012 475322 352064 475328
rect 351920 456000 351972 456006
rect 351920 455942 351972 455948
rect 351552 450832 351604 450838
rect 351552 450774 351604 450780
rect 350920 449942 351210 449970
rect 351564 449956 351592 450774
rect 352024 449970 352052 475322
rect 352746 459776 352802 459785
rect 352746 459711 352802 459720
rect 352380 456000 352432 456006
rect 352380 455942 352432 455948
rect 352286 452024 352342 452033
rect 352286 451959 352342 451968
rect 351946 449942 352052 449970
rect 352300 449956 352328 451959
rect 352392 449970 352420 455942
rect 352760 449970 352788 459711
rect 353312 457842 353340 489126
rect 353392 472796 353444 472802
rect 353392 472738 353444 472744
rect 353300 457836 353352 457842
rect 353300 457778 353352 457784
rect 352392 449942 352682 449970
rect 352760 449942 353050 449970
rect 353404 449956 353432 472738
rect 353852 457836 353904 457842
rect 353852 457778 353904 457784
rect 353760 450424 353812 450430
rect 353760 450366 353812 450372
rect 353772 449956 353800 450366
rect 353864 449970 353892 457778
rect 354692 456006 354720 495406
rect 354772 493400 354824 493406
rect 354772 493342 354824 493348
rect 354680 456000 354732 456006
rect 354680 455942 354732 455948
rect 354494 450120 354550 450129
rect 354494 450055 354550 450064
rect 353864 449942 354154 449970
rect 354508 449956 354536 450055
rect 354784 449970 354812 493342
rect 356060 485240 356112 485246
rect 356060 485182 356112 485188
rect 355690 458688 355746 458697
rect 355690 458623 355746 458632
rect 355324 456000 355376 456006
rect 355324 455942 355376 455948
rect 354956 454368 355008 454374
rect 354956 454310 355008 454316
rect 354968 449970 354996 454310
rect 355336 449970 355364 455942
rect 355704 449970 355732 458623
rect 356072 449970 356100 485182
rect 356152 475380 356204 475386
rect 356152 475322 356204 475328
rect 356164 460934 356192 475322
rect 356164 460906 356836 460934
rect 356704 450560 356756 450566
rect 356704 450502 356756 450508
rect 354784 449942 354890 449970
rect 354968 449942 355258 449970
rect 355336 449942 355626 449970
rect 355704 449942 355994 449970
rect 356072 449942 356362 449970
rect 356716 449956 356744 450502
rect 356808 449970 356836 460906
rect 357452 456006 357480 500142
rect 364076 500138 364104 500686
rect 364616 500686 364668 500692
rect 366362 500712 366418 500721
rect 364154 500647 364210 500656
rect 364064 500132 364116 500138
rect 364064 500074 364116 500080
rect 364628 500070 364656 500686
rect 366362 500647 366418 500656
rect 364616 500064 364668 500070
rect 364616 500006 364668 500012
rect 360476 497412 360528 497418
rect 360476 497354 360528 497360
rect 360292 494896 360344 494902
rect 360292 494838 360344 494844
rect 357532 478304 357584 478310
rect 357532 478246 357584 478252
rect 357440 456000 357492 456006
rect 357440 455942 357492 455948
rect 357438 450256 357494 450265
rect 357438 450191 357494 450200
rect 356808 449942 357098 449970
rect 357452 449956 357480 450191
rect 357544 449970 357572 478246
rect 358820 472660 358872 472666
rect 358820 472602 358872 472608
rect 358832 460934 358860 472602
rect 358832 460906 359780 460934
rect 358912 460284 358964 460290
rect 358912 460226 358964 460232
rect 358268 456000 358320 456006
rect 358268 455942 358320 455948
rect 357900 454844 357952 454850
rect 357900 454786 357952 454792
rect 357912 449970 357940 454786
rect 358280 449970 358308 455942
rect 358924 450498 358952 460226
rect 359002 459640 359058 459649
rect 359002 459575 359058 459584
rect 358912 450492 358964 450498
rect 358912 450434 358964 450440
rect 359016 449970 359044 459575
rect 359648 450560 359700 450566
rect 359648 450502 359700 450508
rect 359096 450492 359148 450498
rect 359096 450434 359148 450440
rect 357544 449942 357834 449970
rect 357912 449942 358202 449970
rect 358280 449942 358570 449970
rect 358938 449942 359044 449970
rect 359108 449970 359136 450434
rect 359108 449942 359306 449970
rect 359660 449956 359688 450502
rect 359752 449970 359780 460906
rect 360200 457088 360252 457094
rect 360200 457030 360252 457036
rect 360212 449970 360240 457030
rect 360304 451274 360332 494838
rect 360488 460934 360516 497354
rect 363236 491972 363288 491978
rect 363236 491914 363288 491920
rect 363052 468512 363104 468518
rect 363052 468454 363104 468460
rect 361580 463208 361632 463214
rect 361580 463150 361632 463156
rect 361592 460934 361620 463150
rect 360488 460906 361252 460934
rect 361592 460906 361988 460934
rect 361120 453484 361172 453490
rect 361120 453426 361172 453432
rect 360304 451246 360516 451274
rect 360488 449970 360516 451246
rect 359752 449942 360042 449970
rect 360212 449942 360410 449970
rect 360488 449942 360778 449970
rect 361132 449956 361160 453426
rect 361224 449970 361252 460906
rect 361670 458552 361726 458561
rect 361670 458487 361726 458496
rect 361684 449970 361712 458487
rect 361960 449970 361988 460906
rect 362592 453416 362644 453422
rect 362592 453358 362644 453364
rect 361224 449942 361514 449970
rect 361684 449942 361882 449970
rect 361960 449942 362250 449970
rect 362604 449956 362632 453358
rect 363064 449970 363092 468454
rect 363248 460934 363276 491914
rect 365904 465792 365956 465798
rect 365904 465734 365956 465740
rect 364340 463140 364392 463146
rect 364340 463082 364392 463088
rect 363248 460906 363460 460934
rect 363144 455864 363196 455870
rect 363144 455806 363196 455812
rect 362986 449942 363092 449970
rect 363156 449970 363184 455806
rect 363432 449970 363460 460906
rect 364352 456006 364380 463082
rect 364430 462496 364486 462505
rect 364430 462431 364486 462440
rect 364444 460934 364472 462431
rect 364444 460906 364564 460934
rect 364340 456000 364392 456006
rect 364340 455942 364392 455948
rect 364432 452260 364484 452266
rect 364432 452202 364484 452208
rect 364062 452160 364118 452169
rect 364062 452095 364118 452104
rect 363156 449942 363354 449970
rect 363432 449942 363722 449970
rect 364076 449956 364104 452095
rect 364444 449956 364472 452202
rect 364536 449970 364564 460906
rect 364892 456000 364944 456006
rect 364892 455942 364944 455948
rect 364904 449970 364932 455942
rect 364536 449942 364826 449970
rect 364904 449942 365194 449970
rect 365562 449954 365760 449970
rect 365916 449956 365944 465734
rect 366376 460934 366404 500647
rect 369122 500032 369178 500041
rect 369122 499967 369178 499976
rect 368756 474088 368808 474094
rect 368756 474030 368808 474036
rect 368572 467152 368624 467158
rect 368572 467094 368624 467100
rect 366284 460906 366404 460934
rect 365996 457020 366048 457026
rect 365996 456962 366048 456968
rect 366008 449970 366036 456962
rect 366284 451994 366312 460906
rect 367836 456204 367888 456210
rect 367836 456146 367888 456152
rect 367468 455048 367520 455054
rect 367468 454990 367520 454996
rect 366364 454708 366416 454714
rect 366364 454650 366416 454656
rect 366272 451988 366324 451994
rect 366272 451930 366324 451936
rect 366376 449970 366404 454650
rect 367376 451988 367428 451994
rect 367376 451930 367428 451936
rect 365562 449948 365772 449954
rect 365562 449942 365720 449948
rect 366008 449942 366298 449970
rect 366376 449942 366666 449970
rect 367388 449956 367416 451930
rect 367480 449970 367508 454990
rect 367848 449970 367876 456146
rect 368480 450628 368532 450634
rect 368480 450570 368532 450576
rect 367480 449942 367770 449970
rect 367848 449942 368138 449970
rect 368492 449956 368520 450570
rect 368584 449970 368612 467094
rect 368768 460934 368796 474030
rect 368768 460906 369072 460934
rect 368940 455796 368992 455802
rect 368940 455738 368992 455744
rect 368756 454912 368808 454918
rect 368756 454854 368808 454860
rect 368768 452169 368796 454854
rect 368754 452160 368810 452169
rect 368754 452095 368810 452104
rect 368952 449970 368980 455738
rect 369044 451274 369072 460906
rect 369136 451926 369164 499967
rect 377600 495106 377628 682042
rect 377680 681896 377732 681902
rect 377680 681838 377732 681844
rect 377692 498030 377720 681838
rect 377784 500041 377812 682654
rect 379704 682644 379756 682650
rect 379704 682586 379756 682592
rect 379612 682508 379664 682514
rect 379612 682450 379664 682456
rect 378324 682440 378376 682446
rect 378324 682382 378376 682388
rect 378232 682304 378284 682310
rect 378232 682246 378284 682252
rect 378138 584760 378194 584769
rect 378138 584695 378194 584704
rect 377862 584488 377918 584497
rect 377862 584423 377918 584432
rect 377770 500032 377826 500041
rect 377770 499967 377826 499976
rect 377680 498024 377732 498030
rect 377680 497966 377732 497972
rect 377588 495100 377640 495106
rect 377588 495042 377640 495048
rect 371240 476876 371292 476882
rect 371240 476818 371292 476824
rect 370134 461136 370190 461145
rect 370134 461071 370190 461080
rect 370148 460934 370176 461071
rect 370148 460906 370452 460934
rect 369860 452600 369912 452606
rect 369860 452542 369912 452548
rect 369872 452062 369900 452542
rect 369950 452432 370006 452441
rect 369950 452367 370006 452376
rect 369860 452056 369912 452062
rect 369860 451998 369912 452004
rect 369124 451920 369176 451926
rect 369124 451862 369176 451868
rect 369044 451246 369348 451274
rect 369320 449970 369348 451246
rect 368584 449942 368874 449970
rect 368952 449942 369242 449970
rect 369320 449942 369610 449970
rect 369964 449956 369992 452367
rect 370320 452260 370372 452266
rect 370320 452202 370372 452208
rect 370332 449956 370360 452202
rect 370424 449970 370452 460906
rect 371056 453620 371108 453626
rect 371056 453562 371108 453568
rect 370424 449942 370714 449970
rect 371068 449956 371096 453562
rect 371252 452674 371280 476818
rect 375380 469940 375432 469946
rect 375380 469882 375432 469888
rect 371332 469872 371384 469878
rect 371332 469814 371384 469820
rect 371344 460934 371372 469814
rect 374000 464432 374052 464438
rect 374000 464374 374052 464380
rect 371344 460906 371556 460934
rect 371240 452668 371292 452674
rect 371240 452610 371292 452616
rect 371424 450696 371476 450702
rect 371424 450638 371476 450644
rect 371436 449956 371464 450638
rect 371528 449970 371556 460906
rect 374012 459542 374040 464374
rect 374092 461780 374144 461786
rect 374092 461722 374144 461728
rect 374000 459536 374052 459542
rect 374000 459478 374052 459484
rect 371882 457192 371938 457201
rect 371882 457127 371938 457136
rect 371896 449970 371924 457127
rect 373630 454608 373686 454617
rect 373630 454543 373686 454552
rect 372252 452668 372304 452674
rect 372252 452610 372304 452616
rect 372264 449970 372292 452610
rect 373262 452568 373318 452577
rect 373262 452503 373318 452512
rect 372434 451888 372490 451897
rect 372434 451823 372490 451832
rect 372448 450809 372476 451823
rect 372528 451716 372580 451722
rect 372528 451658 372580 451664
rect 372896 451716 372948 451722
rect 372896 451658 372948 451664
rect 372434 450800 372490 450809
rect 372434 450735 372490 450744
rect 372540 450673 372568 451658
rect 372526 450664 372582 450673
rect 372526 450599 372582 450608
rect 371528 449942 371818 449970
rect 371896 449942 372186 449970
rect 372264 449942 372554 449970
rect 372908 449956 372936 451658
rect 373276 449956 373304 452503
rect 373644 449956 373672 454543
rect 374104 449970 374132 461722
rect 374460 459536 374512 459542
rect 374460 459478 374512 459484
rect 374368 450764 374420 450770
rect 374368 450706 374420 450712
rect 374026 449942 374132 449970
rect 374380 449956 374408 450706
rect 374472 449970 374500 459478
rect 375102 455832 375158 455841
rect 375102 455767 375158 455776
rect 374472 449942 374762 449970
rect 375116 449956 375144 455767
rect 375392 449970 375420 469882
rect 376760 463072 376812 463078
rect 376760 463014 376812 463020
rect 375470 461000 375526 461009
rect 375470 460935 375526 460944
rect 375484 456794 375512 460935
rect 375484 456766 376340 456794
rect 376206 452568 376262 452577
rect 376206 452503 376262 452512
rect 375838 452296 375894 452305
rect 375838 452231 375894 452240
rect 375392 449942 375498 449970
rect 375852 449956 375880 452231
rect 376220 449956 376248 452503
rect 376312 449970 376340 456766
rect 376772 452674 376800 463014
rect 376850 461680 376906 461689
rect 376850 461615 376906 461624
rect 376760 452668 376812 452674
rect 376760 452610 376812 452616
rect 376864 449970 376892 461615
rect 377770 457056 377826 457065
rect 377770 456991 377826 457000
rect 377404 452668 377456 452674
rect 377404 452610 377456 452616
rect 377312 452396 377364 452402
rect 377312 452338 377364 452344
rect 376312 449942 376602 449970
rect 376864 449942 376970 449970
rect 377324 449956 377352 452338
rect 377416 449970 377444 452610
rect 377784 449970 377812 456991
rect 377876 452198 377904 584423
rect 378152 452674 378180 584695
rect 378244 497690 378272 682246
rect 378336 497758 378364 682382
rect 378508 682372 378560 682378
rect 378508 682314 378560 682320
rect 378416 681828 378468 681834
rect 378416 681770 378468 681776
rect 378428 497826 378456 681770
rect 378520 498098 378548 682314
rect 379520 682032 379572 682038
rect 379520 681974 379572 681980
rect 378796 586214 379100 586242
rect 378508 498092 378560 498098
rect 378508 498034 378560 498040
rect 378416 497820 378468 497826
rect 378416 497762 378468 497768
rect 378324 497752 378376 497758
rect 378324 497694 378376 497700
rect 378232 497684 378284 497690
rect 378232 497626 378284 497632
rect 378232 463004 378284 463010
rect 378232 462946 378284 462952
rect 378140 452668 378192 452674
rect 378140 452610 378192 452616
rect 377864 452192 377916 452198
rect 377864 452134 377916 452140
rect 378138 452024 378194 452033
rect 378138 451959 378194 451968
rect 378152 451858 378180 451959
rect 378140 451852 378192 451858
rect 378140 451794 378192 451800
rect 378244 449970 378272 462946
rect 378796 460934 378824 586214
rect 378704 460906 378824 460934
rect 378888 586090 379008 586106
rect 379072 586090 379100 586214
rect 378888 586084 379020 586090
rect 378888 586078 378968 586084
rect 378704 452606 378732 460906
rect 378888 456794 378916 586078
rect 378968 586026 379020 586032
rect 379060 586084 379112 586090
rect 379060 586026 379112 586032
rect 378968 585948 379020 585954
rect 378968 585890 379020 585896
rect 378796 456766 378916 456794
rect 378692 452600 378744 452606
rect 378692 452542 378744 452548
rect 378796 452130 378824 456766
rect 378876 452668 378928 452674
rect 378876 452610 378928 452616
rect 378784 452124 378836 452130
rect 378784 452066 378836 452072
rect 378782 451888 378838 451897
rect 378782 451823 378838 451832
rect 377416 449942 377706 449970
rect 377784 449942 378074 449970
rect 378244 449942 378442 449970
rect 378796 449956 378824 451823
rect 378888 449970 378916 452610
rect 378980 452266 379008 585890
rect 379060 585812 379112 585818
rect 379060 585754 379112 585760
rect 379072 584769 379100 585754
rect 379058 584760 379114 584769
rect 379058 584695 379114 584704
rect 379058 584624 379114 584633
rect 379058 584559 379114 584568
rect 378968 452260 379020 452266
rect 378968 452202 379020 452208
rect 379072 452062 379100 584559
rect 379152 584452 379204 584458
rect 379152 584394 379204 584400
rect 379060 452056 379112 452062
rect 379060 451998 379112 452004
rect 379164 451926 379192 584394
rect 379532 495038 379560 681974
rect 379624 497894 379652 682450
rect 379612 497888 379664 497894
rect 379612 497830 379664 497836
rect 379716 497554 379744 682586
rect 381176 682576 381228 682582
rect 381176 682518 381228 682524
rect 381084 682236 381136 682242
rect 381084 682178 381136 682184
rect 380992 682168 381044 682174
rect 380992 682110 381044 682116
rect 379796 679040 379848 679046
rect 379796 678982 379848 678988
rect 379808 497962 379836 678982
rect 380164 586560 380216 586566
rect 380164 586502 380216 586508
rect 379796 497956 379848 497962
rect 379796 497898 379848 497904
rect 379704 497548 379756 497554
rect 379704 497490 379756 497496
rect 379520 495032 379572 495038
rect 379520 494974 379572 494980
rect 379520 474088 379572 474094
rect 379520 474030 379572 474036
rect 379532 456210 379560 474030
rect 379610 462360 379666 462369
rect 379610 462295 379666 462304
rect 379520 456204 379572 456210
rect 379520 456146 379572 456152
rect 379152 451920 379204 451926
rect 379152 451862 379204 451868
rect 379624 449970 379652 462295
rect 380176 461718 380204 586502
rect 380900 584520 380952 584526
rect 380900 584462 380952 584468
rect 380164 461712 380216 461718
rect 380164 461654 380216 461660
rect 379702 461544 379758 461553
rect 379702 461479 379758 461488
rect 378888 449942 379178 449970
rect 379546 449942 379652 449970
rect 379716 449970 379744 461479
rect 380912 456210 380940 584462
rect 381004 494970 381032 682110
rect 381096 495174 381124 682178
rect 381188 497622 381216 682518
rect 381268 681964 381320 681970
rect 381268 681906 381320 681912
rect 381280 498982 381308 681906
rect 381268 498976 381320 498982
rect 381268 498918 381320 498924
rect 381176 497616 381228 497622
rect 381176 497558 381228 497564
rect 381084 495168 381136 495174
rect 381084 495110 381136 495116
rect 380992 494964 381044 494970
rect 380992 494906 381044 494912
rect 382936 492114 382964 696934
rect 385684 683188 385736 683194
rect 385684 683130 385736 683136
rect 385040 585880 385092 585886
rect 385040 585822 385092 585828
rect 383016 536104 383068 536110
rect 383016 536046 383068 536052
rect 382924 492108 382976 492114
rect 382924 492050 382976 492056
rect 380992 464364 381044 464370
rect 380992 464306 381044 464312
rect 381004 460934 381032 464306
rect 383028 463690 383056 536046
rect 383660 465724 383712 465730
rect 383660 465666 383712 465672
rect 383016 463684 383068 463690
rect 383016 463626 383068 463632
rect 383672 460934 383700 465666
rect 381004 460906 381216 460934
rect 383672 460906 384068 460934
rect 381084 459604 381136 459610
rect 381084 459546 381136 459552
rect 380348 456204 380400 456210
rect 380348 456146 380400 456152
rect 380900 456204 380952 456210
rect 380900 456146 380952 456152
rect 380256 451920 380308 451926
rect 380256 451862 380308 451868
rect 379716 449942 379914 449970
rect 380268 449956 380296 451862
rect 380360 449970 380388 456146
rect 381096 449970 381124 459546
rect 380360 449942 380650 449970
rect 381018 449942 381124 449970
rect 381188 449970 381216 460906
rect 382554 460184 382610 460193
rect 382554 460119 382610 460128
rect 381820 456204 381872 456210
rect 381820 456146 381872 456152
rect 381728 451308 381780 451314
rect 381728 451250 381780 451256
rect 381188 449942 381386 449970
rect 381740 449956 381768 451250
rect 381832 449970 381860 456146
rect 382370 454472 382426 454481
rect 382370 454407 382426 454416
rect 382384 449970 382412 454407
rect 382568 449970 382596 460119
rect 383292 454708 383344 454714
rect 383292 454650 383344 454656
rect 383200 451512 383252 451518
rect 383200 451454 383252 451460
rect 381832 449942 382122 449970
rect 382384 449942 382490 449970
rect 382568 449942 382858 449970
rect 383212 449956 383240 451454
rect 383304 449970 383332 454650
rect 383660 451376 383712 451382
rect 383660 451318 383712 451324
rect 383672 450945 383700 451318
rect 383658 450936 383714 450945
rect 383658 450871 383714 450880
rect 384040 449970 384068 460906
rect 384672 451376 384724 451382
rect 384672 451318 384724 451324
rect 383304 449942 383594 449970
rect 384040 449942 384330 449970
rect 384684 449956 384712 451318
rect 385052 449956 385080 585822
rect 385696 490822 385724 683130
rect 389178 682136 389234 682145
rect 389178 682071 389234 682080
rect 388166 682000 388222 682009
rect 388166 681935 388222 681944
rect 387064 509924 387116 509930
rect 387064 509866 387116 509872
rect 385776 498840 385828 498846
rect 385776 498782 385828 498788
rect 385684 490816 385736 490822
rect 385684 490758 385736 490764
rect 385130 465760 385186 465769
rect 385130 465695 385186 465704
rect 385144 460934 385172 465695
rect 385144 460906 385540 460934
rect 385408 451308 385460 451314
rect 385408 451250 385460 451256
rect 385420 449956 385448 451250
rect 385512 449970 385540 460906
rect 385788 460902 385816 498782
rect 387076 460902 387104 509866
rect 385776 460896 385828 460902
rect 385776 460838 385828 460844
rect 387064 460896 387116 460902
rect 387064 460838 387116 460844
rect 387076 456210 387104 460838
rect 386144 456204 386196 456210
rect 386144 456146 386196 456152
rect 387064 456204 387116 456210
rect 387064 456146 387116 456152
rect 386156 452674 386184 456146
rect 386144 452668 386196 452674
rect 386144 452610 386196 452616
rect 385512 449942 385802 449970
rect 386156 449956 386184 452610
rect 387616 452532 387668 452538
rect 387616 452474 387668 452480
rect 365720 449890 365772 449896
rect 285706 449806 285996 449834
rect 302266 449806 302556 449834
rect 324346 449806 324636 449834
rect 367006 449848 367062 449857
rect 230478 449783 230534 449792
rect 367006 449783 367062 449792
rect 349620 449744 349672 449750
rect 261390 449712 261446 449721
rect 263520 449682 263626 449698
rect 261390 449647 261446 449656
rect 263508 449676 263626 449682
rect 263560 449670 263626 449676
rect 312570 449682 312860 449698
rect 349370 449692 349620 449698
rect 349370 449686 349672 449692
rect 383934 449712 383990 449721
rect 312570 449676 312872 449682
rect 312570 449670 312820 449676
rect 263508 449618 263560 449624
rect 349370 449670 349660 449686
rect 383934 449647 383990 449656
rect 312820 449618 312872 449624
rect 267464 449608 267516 449614
rect 268568 449608 268620 449614
rect 267516 449556 267674 449562
rect 267464 449550 267674 449556
rect 309048 449608 309100 449614
rect 268620 449556 268778 449562
rect 268568 449550 268778 449556
rect 267476 449534 267674 449550
rect 268580 449534 268778 449550
rect 308890 449556 309048 449562
rect 387628 449585 387656 452474
rect 387708 451648 387760 451654
rect 387708 451590 387760 451596
rect 387720 449818 387748 451590
rect 388076 451308 388128 451314
rect 388076 451250 388128 451256
rect 387708 449812 387760 449818
rect 387708 449754 387760 449760
rect 308890 449550 309100 449556
rect 387614 449576 387670 449585
rect 308890 449534 309088 449550
rect 387614 449511 387670 449520
rect 194046 449304 194102 449313
rect 194046 449239 194102 449248
rect 191838 422376 191894 422385
rect 191838 422311 191894 422320
rect 191838 419656 191894 419665
rect 191838 419591 191894 419600
rect 191852 397361 191880 419591
rect 191838 397352 191894 397361
rect 191838 397287 191894 397296
rect 191838 395992 191894 396001
rect 191838 395927 191894 395936
rect 191852 369209 191880 395927
rect 191838 369200 191894 369209
rect 191838 369135 191894 369144
rect 191838 369064 191894 369073
rect 191838 368999 191894 369008
rect 191748 19032 191800 19038
rect 191748 18974 191800 18980
rect 191656 18760 191708 18766
rect 191656 18702 191708 18708
rect 191472 17808 191524 17814
rect 191472 17750 191524 17756
rect 191852 17610 191880 368999
rect 218704 250504 218756 250510
rect 218704 250446 218756 250452
rect 191944 247722 191972 250036
rect 193324 247790 193352 250036
rect 194612 250022 194718 250050
rect 193312 247784 193364 247790
rect 193312 247726 193364 247732
rect 191932 247716 191984 247722
rect 191932 247658 191984 247664
rect 191840 17604 191892 17610
rect 191840 17546 191892 17552
rect 191378 17504 191434 17513
rect 191378 17439 191434 17448
rect 191104 17060 191156 17066
rect 191104 17002 191156 17008
rect 183572 16546 183784 16574
rect 186332 16546 186912 16574
rect 182916 3664 182968 3670
rect 182916 3606 182968 3612
rect 181352 3596 181404 3602
rect 181352 3538 181404 3544
rect 183756 480 183784 16546
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 194612 4826 194640 250022
rect 196084 247110 196112 250036
rect 197358 247752 197414 247761
rect 197358 247687 197414 247696
rect 195244 247104 195296 247110
rect 195244 247046 195296 247052
rect 196072 247104 196124 247110
rect 196072 247046 196124 247052
rect 195256 10334 195284 247046
rect 195244 10328 195296 10334
rect 195244 10270 195296 10276
rect 197372 6914 197400 247687
rect 197464 14482 197492 250036
rect 198752 250022 198858 250050
rect 198752 15910 198780 250022
rect 200224 248062 200252 250036
rect 201604 248130 201632 250036
rect 202892 250022 202998 250050
rect 201682 248296 201738 248305
rect 201682 248231 201738 248240
rect 201592 248124 201644 248130
rect 201592 248066 201644 248072
rect 200212 248056 200264 248062
rect 200212 247998 200264 248004
rect 201696 238754 201724 248231
rect 201604 238726 201724 238754
rect 198740 15904 198792 15910
rect 198740 15846 198792 15852
rect 197452 14476 197504 14482
rect 197452 14418 197504 14424
rect 201604 6914 201632 238726
rect 197372 6886 197952 6914
rect 194600 4820 194652 4826
rect 194600 4762 194652 4768
rect 194416 3664 194468 3670
rect 194416 3606 194468 3612
rect 190828 3596 190880 3602
rect 190828 3538 190880 3544
rect 190840 480 190868 3538
rect 194428 480 194456 3606
rect 197924 480 197952 6886
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202892 3466 202920 250022
rect 204364 247994 204392 250036
rect 205652 250022 205758 250050
rect 204352 247988 204404 247994
rect 204352 247930 204404 247936
rect 205652 3534 205680 250022
rect 207124 247926 207152 250036
rect 207112 247920 207164 247926
rect 207112 247862 207164 247868
rect 208504 247858 208532 250036
rect 209792 250022 209898 250050
rect 211172 250022 211278 250050
rect 208492 247852 208544 247858
rect 208492 247794 208544 247800
rect 208398 247480 208454 247489
rect 208398 247415 208454 247424
rect 208412 16574 208440 247415
rect 208412 16546 208624 16574
rect 205640 3528 205692 3534
rect 205640 3470 205692 3476
rect 202880 3460 202932 3466
rect 202880 3402 202932 3408
rect 205088 3460 205140 3466
rect 205088 3402 205140 3408
rect 205100 480 205128 3402
rect 208596 480 208624 16546
rect 209792 7614 209820 250022
rect 211172 244934 211200 250022
rect 211252 247648 211304 247654
rect 211252 247590 211304 247596
rect 211160 244928 211212 244934
rect 211160 244870 211212 244876
rect 211264 16574 211292 247590
rect 212644 246362 212672 250036
rect 213932 250022 214038 250050
rect 213182 247888 213238 247897
rect 213182 247823 213238 247832
rect 212632 246356 212684 246362
rect 212632 246298 212684 246304
rect 211264 16546 211752 16574
rect 209780 7608 209832 7614
rect 209780 7550 209832 7556
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213196 3602 213224 247823
rect 213932 6186 213960 250022
rect 214562 248024 214618 248033
rect 214562 247959 214618 247968
rect 213920 6180 213972 6186
rect 213920 6122 213972 6128
rect 214576 3670 214604 247959
rect 215208 247784 215260 247790
rect 215208 247726 215260 247732
rect 215220 3806 215248 247726
rect 215300 247512 215352 247518
rect 215300 247454 215352 247460
rect 215208 3800 215260 3806
rect 215208 3742 215260 3748
rect 214564 3664 214616 3670
rect 214564 3606 214616 3612
rect 213184 3596 213236 3602
rect 213184 3538 213236 3544
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 247454
rect 215404 243574 215432 250036
rect 216404 248396 216456 248402
rect 216404 248338 216456 248344
rect 215942 247344 215998 247353
rect 215942 247279 215998 247288
rect 215392 243568 215444 243574
rect 215392 243510 215444 243516
rect 215956 3466 215984 247279
rect 216220 105732 216272 105738
rect 216220 105674 216272 105680
rect 216128 103556 216180 103562
rect 216128 103498 216180 103504
rect 216140 57934 216168 103498
rect 216128 57928 216180 57934
rect 216128 57870 216180 57876
rect 216232 6390 216260 105674
rect 216312 105664 216364 105670
rect 216312 105606 216364 105612
rect 216220 6384 216272 6390
rect 216220 6326 216272 6332
rect 216324 6254 216352 105606
rect 216312 6248 216364 6254
rect 216312 6190 216364 6196
rect 215944 3460 215996 3466
rect 215944 3402 215996 3408
rect 216416 3262 216444 248338
rect 216588 247852 216640 247858
rect 216588 247794 216640 247800
rect 216496 247716 216548 247722
rect 216496 247658 216548 247664
rect 216508 3670 216536 247658
rect 216600 3738 216628 247794
rect 216784 242214 216812 250036
rect 218072 250022 218178 250050
rect 217322 249112 217378 249121
rect 217322 249047 217378 249056
rect 216772 242208 216824 242214
rect 216772 242150 216824 242156
rect 217232 105800 217284 105806
rect 217232 105742 217284 105748
rect 217140 104236 217192 104242
rect 217140 104178 217192 104184
rect 216680 57928 216732 57934
rect 216680 57870 216732 57876
rect 216692 56953 216720 57870
rect 216678 56944 216734 56953
rect 216678 56879 216734 56888
rect 216680 56568 216732 56574
rect 216680 56510 216732 56516
rect 216692 56001 216720 56510
rect 216678 55992 216734 56001
rect 216678 55927 216734 55936
rect 216678 53816 216734 53825
rect 216678 53751 216680 53760
rect 216732 53751 216734 53760
rect 216680 53722 216732 53728
rect 216772 53712 216824 53718
rect 216772 53654 216824 53660
rect 216784 52873 216812 53654
rect 216770 52864 216826 52873
rect 216770 52799 216826 52808
rect 216772 52420 216824 52426
rect 216772 52362 216824 52368
rect 216784 51105 216812 52362
rect 216770 51096 216826 51105
rect 216680 51060 216732 51066
rect 216770 51031 216826 51040
rect 216680 51002 216732 51008
rect 216692 50017 216720 51002
rect 216678 50008 216734 50017
rect 216678 49943 216734 49952
rect 216680 48272 216732 48278
rect 216678 48240 216680 48249
rect 216732 48240 216734 48249
rect 216678 48175 216734 48184
rect 216588 3732 216640 3738
rect 216588 3674 216640 3680
rect 216496 3664 216548 3670
rect 217152 3641 217180 104178
rect 216496 3606 216548 3612
rect 217138 3632 217194 3641
rect 217138 3567 217194 3576
rect 217244 3505 217272 105742
rect 217336 28529 217364 249047
rect 217600 248328 217652 248334
rect 217600 248270 217652 248276
rect 217508 248260 217560 248266
rect 217508 248202 217560 248208
rect 217416 247580 217468 247586
rect 217416 247522 217468 247528
rect 217322 28520 217378 28529
rect 217322 28455 217378 28464
rect 217322 28384 217378 28393
rect 217322 28319 217378 28328
rect 217336 20058 217364 28319
rect 217324 20052 217376 20058
rect 217324 19994 217376 20000
rect 217428 18426 217456 247522
rect 217416 18420 217468 18426
rect 217416 18362 217468 18368
rect 217230 3496 217286 3505
rect 217230 3431 217286 3440
rect 217520 3398 217548 248202
rect 217508 3392 217560 3398
rect 217508 3334 217560 3340
rect 217612 3330 217640 248270
rect 217968 248192 218020 248198
rect 217968 248134 218020 248140
rect 217876 248124 217928 248130
rect 217876 248066 217928 248072
rect 217784 248056 217836 248062
rect 217784 247998 217836 248004
rect 217692 247920 217744 247926
rect 217692 247862 217744 247868
rect 217704 3942 217732 247862
rect 217796 4010 217824 247998
rect 217888 4078 217916 248066
rect 217980 4146 218008 248134
rect 218072 239426 218100 250022
rect 218060 239420 218112 239426
rect 218060 239362 218112 239368
rect 218060 104168 218112 104174
rect 218060 104110 218112 104116
rect 218072 7614 218100 104110
rect 218716 17134 218744 250446
rect 219452 250022 219558 250050
rect 219348 247988 219400 247994
rect 219348 247930 219400 247936
rect 219164 106004 219216 106010
rect 219164 105946 219216 105952
rect 218980 105596 219032 105602
rect 218980 105538 219032 105544
rect 218704 17128 218756 17134
rect 218704 17070 218756 17076
rect 218888 8356 218940 8362
rect 218888 8298 218940 8304
rect 218060 7608 218112 7614
rect 218060 7550 218112 7556
rect 217968 4140 218020 4146
rect 217968 4082 218020 4088
rect 217876 4072 217928 4078
rect 217876 4014 217928 4020
rect 217784 4004 217836 4010
rect 217784 3946 217836 3952
rect 217692 3936 217744 3942
rect 217692 3878 217744 3884
rect 218900 3369 218928 8298
rect 218992 6186 219020 105538
rect 219072 104372 219124 104378
rect 219072 104314 219124 104320
rect 219084 8362 219112 104314
rect 219072 8356 219124 8362
rect 219072 8298 219124 8304
rect 219176 8242 219204 105946
rect 219256 105868 219308 105874
rect 219256 105810 219308 105816
rect 219084 8214 219204 8242
rect 218980 6180 219032 6186
rect 218980 6122 219032 6128
rect 219084 3602 219112 8214
rect 219268 8106 219296 105810
rect 219176 8078 219296 8106
rect 219176 3913 219204 8078
rect 219256 7608 219308 7614
rect 219256 7550 219308 7556
rect 219162 3904 219218 3913
rect 219162 3839 219218 3848
rect 219072 3596 219124 3602
rect 219072 3538 219124 3544
rect 218886 3360 218942 3369
rect 217600 3324 217652 3330
rect 218886 3295 218942 3304
rect 217600 3266 217652 3272
rect 216404 3256 216456 3262
rect 216404 3198 216456 3204
rect 219268 480 219296 7550
rect 219360 3874 219388 247930
rect 219452 102814 219480 250022
rect 220924 247625 220952 250036
rect 222304 247897 222332 250036
rect 222842 248160 222898 248169
rect 222842 248095 222898 248104
rect 222290 247888 222346 247897
rect 222290 247823 222346 247832
rect 220910 247616 220966 247625
rect 220910 247551 220966 247560
rect 219992 105936 220044 105942
rect 219992 105878 220044 105884
rect 219900 104780 219952 104786
rect 219900 104722 219952 104728
rect 219716 104712 219768 104718
rect 219716 104654 219768 104660
rect 219440 102808 219492 102814
rect 219440 102750 219492 102756
rect 219728 6322 219756 104654
rect 219808 104508 219860 104514
rect 219808 104450 219860 104456
rect 219716 6316 219768 6322
rect 219716 6258 219768 6264
rect 219348 3868 219400 3874
rect 219348 3810 219400 3816
rect 219820 3777 219848 104450
rect 219806 3768 219862 3777
rect 219806 3703 219862 3712
rect 219912 3466 219940 104722
rect 220004 3534 220032 105878
rect 222856 104786 222884 248095
rect 223684 248033 223712 250036
rect 223670 248024 223726 248033
rect 223670 247959 223726 247968
rect 223026 247888 223082 247897
rect 223026 247823 223082 247832
rect 222844 104780 222896 104786
rect 222844 104722 222896 104728
rect 223040 104514 223068 247823
rect 225064 247761 225092 250036
rect 226444 248305 226472 250036
rect 226430 248296 226486 248305
rect 226430 248231 226486 248240
rect 225786 248024 225842 248033
rect 225786 247959 225842 247968
rect 225050 247752 225106 247761
rect 225050 247687 225106 247696
rect 225602 247752 225658 247761
rect 225602 247687 225658 247696
rect 223028 104508 223080 104514
rect 223028 104450 223080 104456
rect 225616 104378 225644 247687
rect 225604 104372 225656 104378
rect 225604 104314 225656 104320
rect 225800 104242 225828 247959
rect 227824 247353 227852 250036
rect 228362 247616 228418 247625
rect 228362 247551 228418 247560
rect 227810 247344 227866 247353
rect 227810 247279 227866 247288
rect 228376 104718 228404 247551
rect 229204 247489 229232 250036
rect 230584 247654 230612 250036
rect 230572 247648 230624 247654
rect 230572 247590 230624 247596
rect 231964 247518 231992 250036
rect 231952 247512 232004 247518
rect 229190 247480 229246 247489
rect 231952 247454 232004 247460
rect 229190 247415 229246 247424
rect 233344 247110 233372 250036
rect 234724 247586 234752 250036
rect 236104 248402 236132 250036
rect 236092 248396 236144 248402
rect 236092 248338 236144 248344
rect 237484 248334 237512 250036
rect 237472 248328 237524 248334
rect 237472 248270 237524 248276
rect 238864 248266 238892 250036
rect 238852 248260 238904 248266
rect 238852 248202 238904 248208
rect 240244 248198 240272 250036
rect 240232 248192 240284 248198
rect 240232 248134 240284 248140
rect 241624 248130 241652 250036
rect 241612 248124 241664 248130
rect 241612 248066 241664 248072
rect 243004 248062 243032 250036
rect 242992 248056 243044 248062
rect 242992 247998 243044 248004
rect 244384 247926 244412 250036
rect 245764 247994 245792 250036
rect 245752 247988 245804 247994
rect 245752 247930 245804 247936
rect 244372 247920 244424 247926
rect 244372 247862 244424 247868
rect 247144 247790 247172 250036
rect 248524 247858 248552 250036
rect 248512 247852 248564 247858
rect 248512 247794 248564 247800
rect 247132 247784 247184 247790
rect 247132 247726 247184 247732
rect 249904 247722 249932 250036
rect 251192 250022 251298 250050
rect 252572 250022 252678 250050
rect 249892 247716 249944 247722
rect 249892 247658 249944 247664
rect 234712 247580 234764 247586
rect 234712 247522 234764 247528
rect 231124 247104 231176 247110
rect 231124 247046 231176 247052
rect 233332 247104 233384 247110
rect 233332 247046 233384 247052
rect 228364 104712 228416 104718
rect 228364 104654 228416 104660
rect 225788 104236 225840 104242
rect 225788 104178 225840 104184
rect 231136 104174 231164 247046
rect 251192 106010 251220 250022
rect 251180 106004 251232 106010
rect 251180 105946 251232 105952
rect 252572 105942 252600 250022
rect 254044 248169 254072 250036
rect 255332 250022 255438 250050
rect 254030 248160 254086 248169
rect 254030 248095 254086 248104
rect 252560 105936 252612 105942
rect 252560 105878 252612 105884
rect 255332 105874 255360 250022
rect 256804 247897 256832 250036
rect 258184 248033 258212 250036
rect 259472 250022 259578 250050
rect 258170 248024 258226 248033
rect 258170 247959 258226 247968
rect 256790 247888 256846 247897
rect 256790 247823 256846 247832
rect 255320 105868 255372 105874
rect 255320 105810 255372 105816
rect 259472 105806 259500 250022
rect 260944 247761 260972 250036
rect 262232 250022 262338 250050
rect 263612 250022 263718 250050
rect 260930 247752 260986 247761
rect 260930 247687 260986 247696
rect 259460 105800 259512 105806
rect 259460 105742 259512 105748
rect 262232 105738 262260 250022
rect 262220 105732 262272 105738
rect 262220 105674 262272 105680
rect 263612 105670 263640 250022
rect 265084 247625 265112 250036
rect 266372 250022 266478 250050
rect 265070 247616 265126 247625
rect 265070 247551 265126 247560
rect 263600 105664 263652 105670
rect 263600 105606 263652 105612
rect 266372 105602 266400 250022
rect 267844 247790 267872 250036
rect 269132 250022 269238 250050
rect 270512 250022 270618 250050
rect 267832 247784 267884 247790
rect 267832 247726 267884 247732
rect 269132 105602 269160 250022
rect 270512 105670 270540 250022
rect 271984 247722 272012 250036
rect 273272 250022 273378 250050
rect 274652 250022 274758 250050
rect 271972 247716 272024 247722
rect 271972 247658 272024 247664
rect 273272 105738 273300 250022
rect 274652 105806 274680 250022
rect 276124 248130 276152 250036
rect 277412 250022 277518 250050
rect 278792 250022 278898 250050
rect 280172 250022 280278 250050
rect 281552 250022 281658 250050
rect 282932 250022 283038 250050
rect 284312 250022 284418 250050
rect 285692 250022 285798 250050
rect 287072 250022 287178 250050
rect 288452 250022 288558 250050
rect 276112 248124 276164 248130
rect 276112 248066 276164 248072
rect 277412 105874 277440 250022
rect 278792 105942 278820 250022
rect 280172 106010 280200 250022
rect 280160 106004 280212 106010
rect 280160 105946 280212 105952
rect 278780 105936 278832 105942
rect 278780 105878 278832 105884
rect 277400 105868 277452 105874
rect 277400 105810 277452 105816
rect 274640 105800 274692 105806
rect 274640 105742 274692 105748
rect 273260 105732 273312 105738
rect 273260 105674 273312 105680
rect 270500 105664 270552 105670
rect 270500 105606 270552 105612
rect 266360 105596 266412 105602
rect 266360 105538 266412 105544
rect 269120 105596 269172 105602
rect 269120 105538 269172 105544
rect 281552 104242 281580 250022
rect 282932 104310 282960 250022
rect 284312 104378 284340 250022
rect 285692 108322 285720 250022
rect 287072 120766 287100 250022
rect 287060 120760 287112 120766
rect 287060 120702 287112 120708
rect 288452 111246 288480 250022
rect 289924 247110 289952 250036
rect 291304 247178 291332 250036
rect 291292 247172 291344 247178
rect 291292 247114 291344 247120
rect 289912 247104 289964 247110
rect 289912 247046 289964 247052
rect 291844 247104 291896 247110
rect 291844 247046 291896 247052
rect 291856 122126 291884 247046
rect 292684 246362 292712 250036
rect 293224 247172 293276 247178
rect 293224 247114 293276 247120
rect 292672 246356 292724 246362
rect 292672 246298 292724 246304
rect 293236 236706 293264 247114
rect 294064 247110 294092 250036
rect 295352 250022 295458 250050
rect 294052 247104 294104 247110
rect 294052 247046 294104 247052
rect 295352 239494 295380 250022
rect 296824 247110 296852 250036
rect 298204 247178 298232 250036
rect 299584 247994 299612 250036
rect 299572 247988 299624 247994
rect 299572 247930 299624 247936
rect 298192 247172 298244 247178
rect 298192 247114 298244 247120
rect 300964 247110 300992 250036
rect 302252 250022 302358 250050
rect 303632 250022 303738 250050
rect 295984 247104 296036 247110
rect 295984 247046 296036 247052
rect 296812 247104 296864 247110
rect 296812 247046 296864 247052
rect 298744 247104 298796 247110
rect 298744 247046 298796 247052
rect 300952 247104 301004 247110
rect 300952 247046 301004 247052
rect 295340 239488 295392 239494
rect 295340 239430 295392 239436
rect 293224 236700 293276 236706
rect 293224 236642 293276 236648
rect 291844 122120 291896 122126
rect 291844 122062 291896 122068
rect 295996 112606 296024 247046
rect 298756 232558 298784 247046
rect 298744 232552 298796 232558
rect 298744 232494 298796 232500
rect 295984 112600 296036 112606
rect 295984 112542 296036 112548
rect 288440 111240 288492 111246
rect 288440 111182 288492 111188
rect 302252 111178 302280 250022
rect 302884 247172 302936 247178
rect 302884 247114 302936 247120
rect 302896 229770 302924 247114
rect 302884 229764 302936 229770
rect 302884 229706 302936 229712
rect 303632 112538 303660 250022
rect 305104 248062 305132 250036
rect 305092 248056 305144 248062
rect 305092 247998 305144 248004
rect 306484 247994 306512 250036
rect 304264 247988 304316 247994
rect 304264 247930 304316 247936
rect 306472 247988 306524 247994
rect 306472 247930 306524 247936
rect 304276 113830 304304 247930
rect 307864 247926 307892 250036
rect 307852 247920 307904 247926
rect 307852 247862 307904 247868
rect 309244 247858 309272 250036
rect 310532 250022 310638 250050
rect 309232 247852 309284 247858
rect 309232 247794 309284 247800
rect 305644 247104 305696 247110
rect 305644 247046 305696 247052
rect 305656 115258 305684 247046
rect 310532 180130 310560 250022
rect 312004 248198 312032 250036
rect 313384 248402 313412 250036
rect 313372 248396 313424 248402
rect 313372 248338 313424 248344
rect 314764 248334 314792 250036
rect 314752 248328 314804 248334
rect 314752 248270 314804 248276
rect 316144 248266 316172 250036
rect 317432 250022 317538 250050
rect 318812 250022 318918 250050
rect 316132 248260 316184 248266
rect 316132 248202 316184 248208
rect 311992 248192 312044 248198
rect 311992 248134 312044 248140
rect 310520 180124 310572 180130
rect 310520 180066 310572 180072
rect 305644 115252 305696 115258
rect 305644 115194 305696 115200
rect 304264 113824 304316 113830
rect 304264 113766 304316 113772
rect 303620 112532 303672 112538
rect 303620 112474 303672 112480
rect 302240 111172 302292 111178
rect 302240 111114 302292 111120
rect 317432 111110 317460 250022
rect 318812 112470 318840 250022
rect 320284 247654 320312 250036
rect 321572 250022 321678 250050
rect 322952 250022 323058 250050
rect 324332 250022 324438 250050
rect 320272 247648 320324 247654
rect 320272 247590 320324 247596
rect 321572 123486 321600 250022
rect 322952 124914 322980 250022
rect 324332 126274 324360 250022
rect 325804 244934 325832 250036
rect 327092 250022 327198 250050
rect 328472 250022 328578 250050
rect 329852 250022 329958 250050
rect 325792 244928 325844 244934
rect 325792 244870 325844 244876
rect 327092 127634 327120 250022
rect 328472 233918 328500 250022
rect 328460 233912 328512 233918
rect 328460 233854 328512 233860
rect 327080 127628 327132 127634
rect 327080 127570 327132 127576
rect 324320 126268 324372 126274
rect 324320 126210 324372 126216
rect 322940 124908 322992 124914
rect 322940 124850 322992 124856
rect 321560 123480 321612 123486
rect 321560 123422 321612 123428
rect 318800 112464 318852 112470
rect 318800 112406 318852 112412
rect 317420 111104 317472 111110
rect 317420 111046 317472 111052
rect 285680 108316 285732 108322
rect 285680 108258 285732 108264
rect 284300 104372 284352 104378
rect 284300 104314 284352 104320
rect 282920 104304 282972 104310
rect 282920 104246 282972 104252
rect 281540 104236 281592 104242
rect 281540 104178 281592 104184
rect 329852 104174 329880 250022
rect 331324 247586 331352 250036
rect 331312 247580 331364 247586
rect 331312 247522 331364 247528
rect 332704 243642 332732 250036
rect 333992 250022 334098 250050
rect 335372 250022 335478 250050
rect 336752 250022 336858 250050
rect 332692 243636 332744 243642
rect 332692 243578 332744 243584
rect 333992 129062 334020 250022
rect 333980 129056 334032 129062
rect 333980 128998 334032 129004
rect 335372 106962 335400 250022
rect 336752 111081 336780 250022
rect 338224 247518 338252 250036
rect 339512 250022 339618 250050
rect 338212 247512 338264 247518
rect 338212 247454 338264 247460
rect 336738 111072 336794 111081
rect 336738 111007 336794 111016
rect 339512 107030 339540 250022
rect 340984 247625 341012 250036
rect 342272 250022 342378 250050
rect 340970 247616 341026 247625
rect 340970 247551 341026 247560
rect 342272 111217 342300 250022
rect 343744 247897 343772 250036
rect 343730 247888 343786 247897
rect 343730 247823 343786 247832
rect 345124 247761 345152 250036
rect 346412 250022 346518 250050
rect 345110 247752 345166 247761
rect 345110 247687 345166 247696
rect 342258 111208 342314 111217
rect 342258 111143 342314 111152
rect 339500 107024 339552 107030
rect 339500 106966 339552 106972
rect 335360 106956 335412 106962
rect 335360 106898 335412 106904
rect 346412 104446 346440 250022
rect 347884 248033 347912 250036
rect 349172 250022 349278 250050
rect 350552 250022 350658 250050
rect 351932 250022 352038 250050
rect 347870 248024 347926 248033
rect 347870 247959 347926 247968
rect 349172 104514 349200 250022
rect 350552 104582 350580 250022
rect 351184 117972 351236 117978
rect 351184 117914 351236 117920
rect 351196 106282 351224 117914
rect 351184 106276 351236 106282
rect 351184 106218 351236 106224
rect 351196 106185 351224 106218
rect 351182 106176 351238 106185
rect 351182 106111 351238 106120
rect 351932 104650 351960 250022
rect 353404 247353 353432 250036
rect 353390 247344 353446 247353
rect 353390 247279 353446 247288
rect 354784 247081 354812 250036
rect 356164 247217 356192 250036
rect 357452 250022 357558 250050
rect 356794 247888 356850 247897
rect 356794 247823 356850 247832
rect 356612 247784 356664 247790
rect 356612 247726 356664 247732
rect 356150 247208 356206 247217
rect 356150 247143 356206 247152
rect 354770 247072 354826 247081
rect 354770 247007 354826 247016
rect 351920 104644 351972 104650
rect 351920 104586 351972 104592
rect 350540 104576 350592 104582
rect 350540 104518 350592 104524
rect 349160 104508 349212 104514
rect 349160 104450 349212 104456
rect 346400 104440 346452 104446
rect 346400 104382 346452 104388
rect 231124 104168 231176 104174
rect 231124 104110 231176 104116
rect 329840 104168 329892 104174
rect 329840 104110 329892 104116
rect 285954 19544 286010 19553
rect 285954 19479 286010 19488
rect 285968 19378 285996 19479
rect 285956 19372 286008 19378
rect 285956 19314 286008 19320
rect 244280 19304 244332 19310
rect 244278 19272 244280 19281
rect 244332 19272 244334 19281
rect 244278 19207 244334 19216
rect 245290 19272 245346 19281
rect 245290 19207 245346 19216
rect 246394 19272 246450 19281
rect 246394 19207 246396 19216
rect 245304 19174 245332 19207
rect 246448 19207 246450 19216
rect 246396 19178 246448 19184
rect 245292 19168 245344 19174
rect 245292 19110 245344 19116
rect 248234 19136 248290 19145
rect 248234 19071 248236 19080
rect 248288 19071 248290 19080
rect 250074 19136 250130 19145
rect 250074 19071 250130 19080
rect 248236 19042 248288 19048
rect 250088 19038 250116 19071
rect 250076 19032 250128 19038
rect 247498 19000 247554 19009
rect 250076 18974 250128 18980
rect 250626 19000 250682 19009
rect 247498 18935 247500 18944
rect 247552 18935 247554 18944
rect 250626 18935 250682 18944
rect 247500 18906 247552 18912
rect 250640 18902 250668 18935
rect 250628 18896 250680 18902
rect 250628 18838 250680 18844
rect 252282 18864 252338 18873
rect 252282 18799 252284 18808
rect 252336 18799 252338 18808
rect 253570 18864 253626 18873
rect 253570 18799 253626 18808
rect 252284 18770 252336 18776
rect 253584 18766 253612 18799
rect 253572 18760 253624 18766
rect 253572 18702 253624 18708
rect 255962 18728 256018 18737
rect 255962 18663 255964 18672
rect 256016 18663 256018 18672
rect 258354 18728 258410 18737
rect 258354 18663 258410 18672
rect 255964 18634 256016 18640
rect 258368 18630 258396 18663
rect 258356 18624 258408 18630
rect 235998 18592 236054 18601
rect 235998 18527 236054 18536
rect 243082 18592 243138 18601
rect 258356 18566 258408 18572
rect 243082 18527 243084 18536
rect 236012 18494 236040 18527
rect 243136 18527 243138 18536
rect 243084 18498 243136 18504
rect 236000 18488 236052 18494
rect 236000 18430 236052 18436
rect 222200 18420 222252 18426
rect 222200 18362 222252 18368
rect 222212 16574 222240 18362
rect 280160 17944 280212 17950
rect 273258 17912 273314 17921
rect 273258 17847 273314 17856
rect 277398 17912 277454 17921
rect 277398 17847 277400 17856
rect 273272 17814 273300 17847
rect 277452 17847 277454 17856
rect 280158 17912 280160 17921
rect 280212 17912 280214 17921
rect 280158 17847 280214 17856
rect 277400 17818 277452 17824
rect 273260 17808 273312 17814
rect 263598 17776 263654 17785
rect 263598 17711 263654 17720
rect 264978 17776 265034 17785
rect 273260 17750 273312 17756
rect 264978 17711 264980 17720
rect 263612 17678 263640 17711
rect 265032 17711 265034 17720
rect 264980 17682 265032 17688
rect 263600 17672 263652 17678
rect 259550 17640 259606 17649
rect 259550 17575 259606 17584
rect 260838 17640 260894 17649
rect 263600 17614 263652 17620
rect 270498 17640 270554 17649
rect 260838 17575 260894 17584
rect 270498 17575 270500 17584
rect 259458 17504 259514 17513
rect 259564 17474 259592 17575
rect 260852 17542 260880 17575
rect 270552 17575 270554 17584
rect 270500 17546 270552 17552
rect 260840 17536 260892 17542
rect 260840 17478 260892 17484
rect 259458 17439 259514 17448
rect 259552 17468 259604 17474
rect 259472 17406 259500 17439
rect 259552 17410 259604 17416
rect 259460 17400 259512 17406
rect 255318 17368 255374 17377
rect 255318 17303 255374 17312
rect 256698 17368 256754 17377
rect 256698 17303 256754 17312
rect 258078 17368 258134 17377
rect 259460 17342 259512 17348
rect 258078 17303 258080 17312
rect 255332 17202 255360 17303
rect 256712 17270 256740 17303
rect 258132 17303 258134 17312
rect 258080 17274 258132 17280
rect 256700 17264 256752 17270
rect 256700 17206 256752 17212
rect 282918 17232 282974 17241
rect 255320 17196 255372 17202
rect 282918 17167 282974 17176
rect 255320 17138 255372 17144
rect 282932 17134 282960 17167
rect 282920 17128 282972 17134
rect 251178 17096 251234 17105
rect 282920 17070 282972 17076
rect 251178 17031 251180 17040
rect 251232 17031 251234 17040
rect 251180 17002 251232 17008
rect 222212 16546 222792 16574
rect 219992 3528 220044 3534
rect 219992 3470 220044 3476
rect 219900 3460 219952 3466
rect 219900 3402 219952 3408
rect 222764 480 222792 16546
rect 293684 6384 293736 6390
rect 293684 6326 293736 6332
rect 237012 4140 237064 4146
rect 237012 4082 237064 4088
rect 233424 3392 233476 3398
rect 233424 3334 233476 3340
rect 229836 3324 229888 3330
rect 229836 3266 229888 3272
rect 226340 3256 226392 3262
rect 226340 3198 226392 3204
rect 226352 480 226380 3198
rect 229848 480 229876 3266
rect 233436 480 233464 3334
rect 237024 480 237052 4082
rect 240508 4072 240560 4078
rect 240508 4014 240560 4020
rect 240520 480 240548 4014
rect 244096 4004 244148 4010
rect 244096 3946 244148 3952
rect 244108 480 244136 3946
rect 247592 3936 247644 3942
rect 247592 3878 247644 3884
rect 276018 3904 276074 3913
rect 247604 480 247632 3878
rect 251180 3868 251232 3874
rect 276018 3839 276074 3848
rect 251180 3810 251232 3816
rect 251192 480 251220 3810
rect 254676 3800 254728 3806
rect 254676 3742 254728 3748
rect 254688 480 254716 3742
rect 258264 3732 258316 3738
rect 258264 3674 258316 3680
rect 258276 480 258304 3674
rect 261760 3664 261812 3670
rect 261760 3606 261812 3612
rect 261772 480 261800 3606
rect 265348 3596 265400 3602
rect 265348 3538 265400 3544
rect 265360 480 265388 3538
rect 268844 3528 268896 3534
rect 268844 3470 268896 3476
rect 268856 480 268884 3470
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 272444 480 272472 3402
rect 276032 480 276060 3839
rect 279514 3768 279570 3777
rect 279514 3703 279570 3712
rect 279528 480 279556 3703
rect 283102 3632 283158 3641
rect 283102 3567 283158 3576
rect 283116 480 283144 3567
rect 286598 3496 286654 3505
rect 286598 3431 286654 3440
rect 286612 480 286640 3431
rect 290186 3360 290242 3369
rect 290186 3295 290242 3304
rect 290200 480 290228 3295
rect 293696 480 293724 6326
rect 300768 6316 300820 6322
rect 300768 6258 300820 6264
rect 297272 6248 297324 6254
rect 297272 6190 297324 6196
rect 297284 480 297312 6190
rect 300780 480 300808 6258
rect 304356 6180 304408 6186
rect 304356 6122 304408 6128
rect 304368 480 304396 6122
rect 343364 4140 343416 4146
rect 343364 4082 343416 4088
rect 339868 4072 339920 4078
rect 339868 4014 339920 4020
rect 336280 4004 336332 4010
rect 336280 3946 336332 3952
rect 332692 3936 332744 3942
rect 332692 3878 332744 3884
rect 329196 3868 329248 3874
rect 329196 3810 329248 3816
rect 325608 3800 325660 3806
rect 325608 3742 325660 3748
rect 322112 3732 322164 3738
rect 322112 3674 322164 3680
rect 318524 3664 318576 3670
rect 318524 3606 318576 3612
rect 315028 3596 315080 3602
rect 315028 3538 315080 3544
rect 311440 3528 311492 3534
rect 311440 3470 311492 3476
rect 307944 3460 307996 3466
rect 307944 3402 307996 3408
rect 307956 480 307984 3402
rect 311452 480 311480 3470
rect 315040 480 315068 3538
rect 318536 480 318564 3606
rect 322124 480 322152 3674
rect 325620 480 325648 3742
rect 329208 480 329236 3810
rect 332704 480 332732 3878
rect 336292 480 336320 3946
rect 339880 480 339908 4014
rect 343376 480 343404 4082
rect 356624 3466 356652 247726
rect 356704 247512 356756 247518
rect 356704 247454 356756 247460
rect 356716 5302 356744 247454
rect 356704 5296 356756 5302
rect 356704 5238 356756 5244
rect 356808 5166 356836 247823
rect 357162 247344 357218 247353
rect 357162 247279 357218 247288
rect 356978 247072 357034 247081
rect 356978 247007 357034 247016
rect 356992 98802 357020 247007
rect 357072 105732 357124 105738
rect 357072 105674 357124 105680
rect 356980 98796 357032 98802
rect 356980 98738 357032 98744
rect 357084 98682 357112 105674
rect 356900 98654 357112 98682
rect 357176 98666 357204 247279
rect 357256 106004 357308 106010
rect 357256 105946 357308 105952
rect 357164 98660 357216 98666
rect 356796 5160 356848 5166
rect 356796 5102 356848 5108
rect 356900 3738 356928 98654
rect 357164 98602 357216 98608
rect 356980 98592 357032 98598
rect 357268 98546 357296 105946
rect 356980 98534 357032 98540
rect 356992 7614 357020 98534
rect 357084 98518 357296 98546
rect 356980 7608 357032 7614
rect 356980 7550 357032 7556
rect 357084 4078 357112 98518
rect 357164 98456 357216 98462
rect 357164 98398 357216 98404
rect 357176 7682 357204 98398
rect 357452 11898 357480 250022
rect 358360 248396 358412 248402
rect 358360 248338 358412 248344
rect 357532 248124 357584 248130
rect 357532 248066 357584 248072
rect 357440 11892 357492 11898
rect 357440 11834 357492 11840
rect 357544 11778 357572 248066
rect 358082 248024 358138 248033
rect 358082 247959 358138 247968
rect 357624 120760 357676 120766
rect 357624 120702 357676 120708
rect 357452 11750 357572 11778
rect 357164 7676 357216 7682
rect 357164 7618 357216 7624
rect 357072 4072 357124 4078
rect 357072 4014 357124 4020
rect 357452 3874 357480 11750
rect 357636 11642 357664 120702
rect 357900 105936 357952 105942
rect 357900 105878 357952 105884
rect 357716 105868 357768 105874
rect 357716 105810 357768 105816
rect 357544 11614 357664 11642
rect 357440 3868 357492 3874
rect 357440 3810 357492 3816
rect 356888 3732 356940 3738
rect 356888 3674 356940 3680
rect 356612 3460 356664 3466
rect 356612 3402 356664 3408
rect 346952 3392 347004 3398
rect 346952 3334 347004 3340
rect 346964 480 346992 3334
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 350460 480 350488 3266
rect 354036 3256 354088 3262
rect 354036 3198 354088 3204
rect 354048 480 354076 3198
rect 357544 480 357572 11614
rect 357624 11552 357676 11558
rect 357624 11494 357676 11500
rect 357636 6186 357664 11494
rect 357624 6180 357676 6186
rect 357624 6122 357676 6128
rect 357728 3942 357756 105810
rect 357808 105800 357860 105806
rect 357808 105742 357860 105748
rect 357716 3936 357768 3942
rect 357716 3878 357768 3884
rect 357820 3806 357848 105742
rect 357912 4010 357940 105878
rect 358096 5030 358124 247959
rect 358266 247752 358322 247761
rect 358266 247687 358322 247696
rect 358176 247648 358228 247654
rect 358176 247590 358228 247596
rect 358188 14482 358216 247590
rect 358176 14476 358228 14482
rect 358176 14418 358228 14424
rect 358280 5098 358308 247687
rect 358372 14550 358400 248338
rect 358924 247081 358952 250036
rect 360212 250022 360318 250050
rect 361592 250022 361698 250050
rect 362972 250022 363078 250050
rect 364352 250022 364458 250050
rect 365732 250022 365838 250050
rect 367112 250022 367218 250050
rect 359556 248192 359608 248198
rect 359556 248134 359608 248140
rect 359464 247580 359516 247586
rect 359464 247522 359516 247528
rect 358910 247072 358966 247081
rect 358910 247007 358966 247016
rect 358820 108316 358872 108322
rect 358820 108258 358872 108264
rect 358360 14544 358412 14550
rect 358360 14486 358412 14492
rect 358268 5092 358320 5098
rect 358268 5034 358320 5040
rect 358084 5024 358136 5030
rect 358084 4966 358136 4972
rect 357900 4004 357952 4010
rect 357900 3946 357952 3952
rect 357808 3800 357860 3806
rect 357808 3742 357860 3748
rect 358832 3262 358860 108258
rect 358912 105664 358964 105670
rect 358912 105606 358964 105612
rect 358924 3602 358952 105606
rect 359004 105596 359056 105602
rect 359004 105538 359056 105544
rect 358912 3596 358964 3602
rect 358912 3538 358964 3544
rect 359016 3534 359044 105538
rect 359096 104372 359148 104378
rect 359096 104314 359148 104320
rect 359004 3528 359056 3534
rect 359004 3470 359056 3476
rect 359108 3330 359136 104314
rect 359280 104304 359332 104310
rect 359280 104246 359332 104252
rect 359188 104236 359240 104242
rect 359188 104178 359240 104184
rect 359200 4146 359228 104178
rect 359188 4140 359240 4146
rect 359188 4082 359240 4088
rect 359292 3398 359320 104246
rect 359476 11762 359504 247522
rect 359568 15978 359596 248134
rect 359648 107024 359700 107030
rect 359648 106966 359700 106972
rect 359556 15972 359608 15978
rect 359556 15914 359608 15920
rect 359464 11756 359516 11762
rect 359464 11698 359516 11704
rect 359660 3466 359688 106966
rect 359740 103556 359792 103562
rect 359740 103498 359792 103504
rect 359752 99249 359780 103498
rect 360108 99340 360160 99346
rect 360108 99282 360160 99288
rect 360120 99249 360148 99282
rect 359738 99240 359794 99249
rect 359738 99175 359794 99184
rect 360106 99240 360162 99249
rect 360106 99175 360162 99184
rect 360212 8974 360240 250022
rect 360936 248328 360988 248334
rect 360936 248270 360988 248276
rect 360842 247616 360898 247625
rect 360842 247551 360898 247560
rect 360292 111240 360344 111246
rect 360292 111182 360344 111188
rect 360304 16574 360332 111182
rect 360304 16546 360792 16574
rect 360200 8968 360252 8974
rect 360200 8910 360252 8916
rect 360764 3482 360792 16546
rect 360856 5234 360884 247551
rect 360948 11830 360976 248270
rect 360936 11824 360988 11830
rect 360936 11766 360988 11772
rect 361592 10334 361620 250022
rect 361672 247716 361724 247722
rect 361672 247658 361724 247664
rect 361580 10328 361632 10334
rect 361580 10270 361632 10276
rect 360844 5228 360896 5234
rect 360844 5170 360896 5176
rect 361684 3670 361712 247658
rect 362972 13122 363000 250022
rect 363604 248260 363656 248266
rect 363604 248202 363656 248208
rect 363616 15910 363644 248202
rect 363604 15904 363656 15910
rect 363604 15846 363656 15852
rect 362960 13116 363012 13122
rect 362960 13058 363012 13064
rect 364352 4962 364380 250022
rect 364432 122120 364484 122126
rect 364432 122062 364484 122068
rect 364444 16574 364472 122062
rect 364444 16546 364656 16574
rect 364340 4956 364392 4962
rect 364340 4898 364392 4904
rect 361672 3664 361724 3670
rect 361672 3606 361724 3612
rect 359648 3460 359700 3466
rect 360764 3454 361160 3482
rect 359648 3402 359700 3408
rect 359280 3392 359332 3398
rect 359280 3334 359332 3340
rect 359096 3324 359148 3330
rect 359096 3266 359148 3272
rect 358820 3256 358872 3262
rect 358820 3198 358872 3204
rect 361132 480 361160 3454
rect 364628 480 364656 16546
rect 365732 4894 365760 250022
rect 365720 4888 365772 4894
rect 365720 4830 365772 4836
rect 367112 4758 367140 250022
rect 368584 243574 368612 250036
rect 369872 250022 369978 250050
rect 368572 243568 368624 243574
rect 368572 243510 368624 243516
rect 367192 236700 367244 236706
rect 367192 236642 367244 236648
rect 367204 16574 367232 236642
rect 369872 198014 369900 250022
rect 371240 246356 371292 246362
rect 371240 246298 371292 246304
rect 369860 198008 369912 198014
rect 369860 197950 369912 197956
rect 371148 28280 371200 28286
rect 371148 28222 371200 28228
rect 371160 20058 371188 28222
rect 371148 20052 371200 20058
rect 371148 19994 371200 20000
rect 367204 16546 367784 16574
rect 367100 4752 367152 4758
rect 367100 4694 367152 4700
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 246298
rect 371344 242214 371372 250036
rect 372632 250022 372738 250050
rect 374012 250022 374118 250050
rect 375392 250022 375498 250050
rect 371332 242208 371384 242214
rect 371332 242150 371384 242156
rect 372632 239426 372660 250022
rect 372620 239420 372672 239426
rect 372620 239362 372672 239368
rect 374012 236706 374040 250022
rect 374000 236700 374052 236706
rect 374000 236642 374052 236648
rect 375392 199442 375420 250022
rect 376864 247722 376892 250036
rect 378244 249762 378272 250036
rect 378232 249756 378284 249762
rect 378232 249698 378284 249704
rect 379624 248198 379652 250036
rect 379612 248192 379664 248198
rect 379612 248134 379664 248140
rect 381004 248130 381032 250036
rect 382384 248266 382412 250036
rect 383764 248402 383792 250036
rect 383752 248396 383804 248402
rect 383752 248338 383804 248344
rect 385144 248334 385172 250036
rect 386420 249756 386472 249762
rect 386420 249698 386472 249704
rect 386432 248470 386460 249698
rect 386420 248464 386472 248470
rect 386420 248406 386472 248412
rect 385132 248328 385184 248334
rect 385132 248270 385184 248276
rect 382372 248260 382424 248266
rect 382372 248202 382424 248208
rect 380992 248124 381044 248130
rect 380992 248066 381044 248072
rect 376852 247716 376904 247722
rect 376852 247658 376904 247664
rect 386432 246362 386460 248406
rect 387904 247790 387932 250036
rect 387892 247784 387944 247790
rect 387892 247726 387944 247732
rect 386420 246356 386472 246362
rect 386420 246298 386472 246304
rect 387904 245682 387932 247726
rect 387064 245676 387116 245682
rect 387064 245618 387116 245624
rect 387892 245676 387944 245682
rect 387892 245618 387944 245624
rect 381544 243636 381596 243642
rect 381544 243578 381596 243584
rect 378140 239488 378192 239494
rect 378140 239430 378192 239436
rect 375380 199436 375432 199442
rect 375380 199378 375432 199384
rect 374000 112600 374052 112606
rect 374000 112542 374052 112548
rect 374012 2786 374040 112542
rect 378152 16574 378180 239430
rect 378152 16546 378456 16574
rect 374000 2780 374052 2786
rect 374000 2722 374052 2728
rect 375288 2780 375340 2786
rect 375288 2722 375340 2728
rect 375300 480 375328 2722
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 381556 3602 381584 243578
rect 382280 232552 382332 232558
rect 382280 232494 382332 232500
rect 382292 16574 382320 232494
rect 385040 229764 385092 229770
rect 385040 229706 385092 229712
rect 385052 16574 385080 229706
rect 387076 99346 387104 245618
rect 387064 99340 387116 99346
rect 387064 99282 387116 99288
rect 388088 16590 388116 451250
rect 388180 248266 388208 681935
rect 388442 587208 388498 587217
rect 388442 587143 388498 587152
rect 388456 467294 388484 587143
rect 388444 467288 388496 467294
rect 388444 467230 388496 467236
rect 388628 451920 388680 451926
rect 388628 451862 388680 451868
rect 388442 450528 388498 450537
rect 388442 450463 388498 450472
rect 388168 248260 388220 248266
rect 388168 248202 388220 248208
rect 388456 17785 388484 450463
rect 388536 449948 388588 449954
rect 388536 449890 388588 449896
rect 388548 106729 388576 449890
rect 388640 108322 388668 451862
rect 388812 451784 388864 451790
rect 388812 451726 388864 451732
rect 388718 449984 388774 449993
rect 388718 449919 388774 449928
rect 388628 108316 388680 108322
rect 388628 108258 388680 108264
rect 388732 107409 388760 449919
rect 388824 109138 388852 451726
rect 388904 451580 388956 451586
rect 388904 451522 388956 451528
rect 388916 442270 388944 451522
rect 388996 449812 389048 449818
rect 388996 449754 389048 449760
rect 389008 449546 389036 449754
rect 388996 449540 389048 449546
rect 388996 449482 389048 449488
rect 388904 442264 388956 442270
rect 388904 442206 388956 442212
rect 389192 248402 389220 682071
rect 389272 681760 389324 681766
rect 389272 681702 389324 681708
rect 389180 248396 389232 248402
rect 389180 248338 389232 248344
rect 389284 248334 389312 681702
rect 389364 498228 389416 498234
rect 389364 498170 389416 498176
rect 389376 248470 389404 498170
rect 389836 496194 389864 700266
rect 390558 681864 390614 681873
rect 390558 681799 390614 681808
rect 389916 507884 389968 507890
rect 389916 507826 389968 507832
rect 389928 499526 389956 507826
rect 389916 499520 389968 499526
rect 389916 499462 389968 499468
rect 389928 498234 389956 499462
rect 389916 498228 389968 498234
rect 389916 498170 389968 498176
rect 389824 496188 389876 496194
rect 389824 496130 389876 496136
rect 390284 454572 390336 454578
rect 390284 454514 390336 454520
rect 390100 452736 390152 452742
rect 390100 452678 390152 452684
rect 389916 451852 389968 451858
rect 389916 451794 389968 451800
rect 389824 451444 389876 451450
rect 389824 451386 389876 451392
rect 389364 248464 389416 248470
rect 389364 248406 389416 248412
rect 389272 248328 389324 248334
rect 389272 248270 389324 248276
rect 389180 113824 389232 113830
rect 389180 113766 389232 113772
rect 388812 109132 388864 109138
rect 388812 109074 388864 109080
rect 388718 107400 388774 107409
rect 388718 107335 388774 107344
rect 388534 106720 388590 106729
rect 388534 106655 388590 106664
rect 388442 17776 388498 17785
rect 388442 17711 388498 17720
rect 388076 16584 388128 16590
rect 382292 16546 382412 16574
rect 385052 16546 386000 16574
rect 381544 3596 381596 3602
rect 381544 3538 381596 3544
rect 382384 480 382412 16546
rect 385972 480 386000 16546
rect 389192 16574 389220 113766
rect 389836 18698 389864 451386
rect 389928 18766 389956 451794
rect 390008 451376 390060 451382
rect 390008 451318 390060 451324
rect 389916 18760 389968 18766
rect 389916 18702 389968 18708
rect 389824 18692 389876 18698
rect 389824 18634 389876 18640
rect 390020 18630 390048 451318
rect 390112 107137 390140 452678
rect 390192 452464 390244 452470
rect 390192 452406 390244 452412
rect 390204 142769 390232 452406
rect 390296 379506 390324 454514
rect 390374 451480 390430 451489
rect 390374 451415 390430 451424
rect 390388 422958 390416 451415
rect 390376 422952 390428 422958
rect 390376 422894 390428 422900
rect 390284 379500 390336 379506
rect 390284 379442 390336 379448
rect 390572 248130 390600 681799
rect 391216 497457 391244 700538
rect 393964 700460 394016 700466
rect 393964 700402 394016 700408
rect 392584 700392 392636 700398
rect 392584 700334 392636 700340
rect 391940 497480 391992 497486
rect 391202 497448 391258 497457
rect 391940 497422 391992 497428
rect 391202 497383 391258 497392
rect 391296 455728 391348 455734
rect 391296 455670 391348 455676
rect 391204 452940 391256 452946
rect 391204 452882 391256 452888
rect 390652 452668 390704 452674
rect 390652 452610 390704 452616
rect 390560 248124 390612 248130
rect 390560 248066 390612 248072
rect 390190 142760 390246 142769
rect 390190 142695 390246 142704
rect 390098 107128 390154 107137
rect 390098 107063 390154 107072
rect 390664 104854 390692 452610
rect 390652 104848 390704 104854
rect 390652 104790 390704 104796
rect 391216 28966 391244 452882
rect 391308 325650 391336 455670
rect 391296 325644 391348 325650
rect 391296 325586 391348 325592
rect 391952 248198 391980 497422
rect 392596 475590 392624 700334
rect 392584 475584 392636 475590
rect 392584 475526 392636 475532
rect 393976 462913 394004 700402
rect 397472 700330 397500 703520
rect 410524 700528 410576 700534
rect 410524 700470 410576 700476
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 400864 700324 400916 700330
rect 400864 700266 400916 700272
rect 393962 462904 394018 462913
rect 393962 462839 394018 462848
rect 399668 458652 399720 458658
rect 399668 458594 399720 458600
rect 399484 458584 399536 458590
rect 399484 458526 399536 458532
rect 394148 456952 394200 456958
rect 394148 456894 394200 456900
rect 392676 454504 392728 454510
rect 392676 454446 392728 454452
rect 392584 452804 392636 452810
rect 392584 452746 392636 452752
rect 391940 248192 391992 248198
rect 391940 248134 391992 248140
rect 391940 115252 391992 115258
rect 391940 115194 391992 115200
rect 391204 28960 391256 28966
rect 391204 28902 391256 28908
rect 390008 18624 390060 18630
rect 390008 18566 390060 18572
rect 391952 16574 391980 115194
rect 392596 107642 392624 452746
rect 392688 245614 392716 454446
rect 394056 454436 394108 454442
rect 394056 454378 394108 454384
rect 393964 453688 394016 453694
rect 393964 453630 394016 453636
rect 392676 245608 392728 245614
rect 392676 245550 392728 245556
rect 392584 107636 392636 107642
rect 392584 107578 392636 107584
rect 393976 17066 394004 453630
rect 394068 206990 394096 454378
rect 394160 419490 394188 456894
rect 395436 455660 395488 455666
rect 395436 455602 395488 455608
rect 395344 455592 395396 455598
rect 395344 455534 395396 455540
rect 394148 419484 394200 419490
rect 394148 419426 394200 419432
rect 395356 273222 395384 455534
rect 395448 353258 395476 455602
rect 396724 455524 396776 455530
rect 396724 455466 396776 455472
rect 395436 353252 395488 353258
rect 395436 353194 395488 353200
rect 395344 273216 395396 273222
rect 395344 273158 395396 273164
rect 396736 259418 396764 455466
rect 396724 259412 396776 259418
rect 396724 259354 396776 259360
rect 394056 206984 394108 206990
rect 394056 206926 394108 206932
rect 398840 112532 398892 112538
rect 398840 112474 398892 112480
rect 396080 111172 396132 111178
rect 396080 111114 396132 111120
rect 393964 17060 394016 17066
rect 393964 17002 394016 17008
rect 389192 16546 389496 16574
rect 391952 16546 392624 16574
rect 388076 16526 388128 16532
rect 389468 480 389496 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 111114
rect 398852 3534 398880 112474
rect 399496 19106 399524 458526
rect 399576 458516 399628 458522
rect 399576 458458 399628 458464
rect 399484 19100 399536 19106
rect 399484 19042 399536 19048
rect 399588 19038 399616 458458
rect 399576 19032 399628 19038
rect 399576 18974 399628 18980
rect 399680 18873 399708 458594
rect 400876 457774 400904 700266
rect 407764 699712 407816 699718
rect 407764 699654 407816 699660
rect 403624 597576 403676 597582
rect 403624 597518 403676 597524
rect 403636 475522 403664 597518
rect 406384 537532 406436 537538
rect 406384 537474 406436 537480
rect 403624 475516 403676 475522
rect 403624 475458 403676 475464
rect 406396 473346 406424 537474
rect 407776 500313 407804 699654
rect 407854 533352 407910 533361
rect 407854 533287 407910 533296
rect 407762 500304 407818 500313
rect 407762 500239 407818 500248
rect 405648 473340 405700 473346
rect 405648 473282 405700 473288
rect 406384 473340 406436 473346
rect 406384 473282 406436 473288
rect 405660 472054 405688 473282
rect 405648 472048 405700 472054
rect 405648 471990 405700 471996
rect 402244 458788 402296 458794
rect 402244 458730 402296 458736
rect 400864 457768 400916 457774
rect 400864 457710 400916 457716
rect 399760 456884 399812 456890
rect 399760 456826 399812 456832
rect 399772 365702 399800 456826
rect 399760 365696 399812 365702
rect 399760 365638 399812 365644
rect 399666 18864 399722 18873
rect 399666 18799 399722 18808
rect 402256 18737 402284 458730
rect 402336 458720 402388 458726
rect 402336 458662 402388 458668
rect 402348 19553 402376 458662
rect 403624 456816 403676 456822
rect 403624 456758 403676 456764
rect 402520 454912 402572 454918
rect 402520 454854 402572 454860
rect 402428 452872 402480 452878
rect 402428 452814 402480 452820
rect 402334 19544 402390 19553
rect 402334 19479 402390 19488
rect 402242 18728 402298 18737
rect 402242 18663 402298 18672
rect 402440 17950 402468 452814
rect 402532 18834 402560 454854
rect 402796 454844 402848 454850
rect 402796 454786 402848 454792
rect 402704 454368 402756 454374
rect 402704 454310 402756 454316
rect 402612 453484 402664 453490
rect 402612 453426 402664 453432
rect 402624 18902 402652 453426
rect 402716 19446 402744 454310
rect 402704 19440 402756 19446
rect 402704 19382 402756 19388
rect 402808 19378 402836 454786
rect 403636 313274 403664 456758
rect 405096 454776 405148 454782
rect 405096 454718 405148 454724
rect 405004 454640 405056 454646
rect 405004 454582 405056 454588
rect 403624 313268 403676 313274
rect 403624 313210 403676 313216
rect 402980 248056 403032 248062
rect 402980 247998 403032 248004
rect 402796 19372 402848 19378
rect 402796 19314 402848 19320
rect 402612 18896 402664 18902
rect 402612 18838 402664 18844
rect 402520 18828 402572 18834
rect 402520 18770 402572 18776
rect 402428 17944 402480 17950
rect 402428 17886 402480 17892
rect 402992 16574 403020 247998
rect 405016 17649 405044 454582
rect 405108 19650 405136 454718
rect 405280 453348 405332 453354
rect 405280 453290 405332 453296
rect 405188 453144 405240 453150
rect 405188 453086 405240 453092
rect 405096 19644 405148 19650
rect 405096 19586 405148 19592
rect 405002 17640 405058 17649
rect 405002 17575 405058 17584
rect 405200 17513 405228 453086
rect 405292 19582 405320 453290
rect 405372 453280 405424 453286
rect 405372 453222 405424 453228
rect 405280 19576 405332 19582
rect 405280 19518 405332 19524
rect 405384 19417 405412 453222
rect 405462 450392 405518 450401
rect 405462 450327 405518 450336
rect 405476 19718 405504 450327
rect 405556 449744 405608 449750
rect 405556 449686 405608 449692
rect 405464 19712 405516 19718
rect 405464 19654 405516 19660
rect 405568 19514 405596 449686
rect 405660 146946 405688 471990
rect 407868 469198 407896 533287
rect 410536 500177 410564 700470
rect 413664 699718 413692 703520
rect 429856 700602 429884 703520
rect 429844 700596 429896 700602
rect 429844 700538 429896 700544
rect 462332 700505 462360 703520
rect 462318 700496 462374 700505
rect 478524 700466 478552 703520
rect 494808 700534 494836 703520
rect 494796 700528 494848 700534
rect 494796 700470 494848 700476
rect 462318 700431 462374 700440
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 543476 700369 543504 703520
rect 527180 700334 527232 700340
rect 543462 700360 543518 700369
rect 559668 700330 559696 703520
rect 543462 700295 543518 700304
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 413652 699712 413704 699718
rect 413652 699654 413704 699660
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 551006 674928 551062 674937
rect 551006 674863 551008 674872
rect 551060 674863 551062 674872
rect 557540 674892 557592 674898
rect 551008 674834 551060 674840
rect 557540 674834 557592 674840
rect 417514 626920 417570 626929
rect 417514 626855 417570 626864
rect 417146 625968 417202 625977
rect 417146 625903 417202 625912
rect 416778 598088 416834 598097
rect 416778 598023 416834 598032
rect 416792 597582 416820 598023
rect 416780 597576 416832 597582
rect 416780 597518 416832 597524
rect 414664 587580 414716 587586
rect 414664 587522 414716 587528
rect 413928 587104 413980 587110
rect 413928 587046 413980 587052
rect 413744 587036 413796 587042
rect 413744 586978 413796 586984
rect 413282 584760 413338 584769
rect 413282 584695 413338 584704
rect 411904 530664 411956 530670
rect 411904 530606 411956 530612
rect 410616 530596 410668 530602
rect 410616 530538 410668 530544
rect 410522 500168 410578 500177
rect 410522 500103 410578 500112
rect 407856 469192 407908 469198
rect 407856 469134 407908 469140
rect 410628 465594 410656 530538
rect 411916 466478 411944 530606
rect 413296 498166 413324 584695
rect 413284 498160 413336 498166
rect 413284 498102 413336 498108
rect 413756 495242 413784 586978
rect 413836 586900 413888 586906
rect 413836 586842 413888 586848
rect 413744 495236 413796 495242
rect 413744 495178 413796 495184
rect 413848 490890 413876 586842
rect 413836 490884 413888 490890
rect 413836 490826 413888 490832
rect 413940 484362 413968 587046
rect 414572 533724 414624 533730
rect 414572 533666 414624 533672
rect 413928 484356 413980 484362
rect 413928 484298 413980 484304
rect 414584 469266 414612 533666
rect 414676 474162 414704 587522
rect 416044 586628 416096 586634
rect 416044 586570 416096 586576
rect 415860 586152 415912 586158
rect 415860 586094 415912 586100
rect 414848 584248 414900 584254
rect 414848 584190 414900 584196
rect 414756 583500 414808 583506
rect 414756 583442 414808 583448
rect 414664 474156 414716 474162
rect 414664 474098 414716 474104
rect 413928 469260 413980 469266
rect 413928 469202 413980 469208
rect 414572 469260 414624 469266
rect 414572 469202 414624 469208
rect 411168 466472 411220 466478
rect 411168 466414 411220 466420
rect 411904 466472 411956 466478
rect 411904 466414 411956 466420
rect 409788 465588 409840 465594
rect 409788 465530 409840 465536
rect 410616 465588 410668 465594
rect 410616 465530 410668 465536
rect 409800 465186 409828 465530
rect 409788 465180 409840 465186
rect 409788 465122 409840 465128
rect 407764 454300 407816 454306
rect 407764 454242 407816 454248
rect 407672 449676 407724 449682
rect 407672 449618 407724 449624
rect 407120 247988 407172 247994
rect 407120 247930 407172 247936
rect 405648 146940 405700 146946
rect 405648 146882 405700 146888
rect 406384 129056 406436 129062
rect 406384 128998 406436 129004
rect 405556 19508 405608 19514
rect 405556 19450 405608 19456
rect 405370 19408 405426 19417
rect 405370 19343 405426 19352
rect 405186 17504 405242 17513
rect 405186 17439 405242 17448
rect 402992 16546 403664 16574
rect 398840 3528 398892 3534
rect 398840 3470 398892 3476
rect 400128 3528 400180 3534
rect 400128 3470 400180 3476
rect 400140 480 400168 3470
rect 403636 480 403664 16546
rect 406396 3670 406424 128998
rect 407132 16574 407160 247930
rect 407684 109177 407712 449618
rect 407670 109168 407726 109177
rect 407670 109103 407726 109112
rect 407776 17377 407804 454242
rect 407948 454232 408000 454238
rect 407948 454174 408000 454180
rect 407856 453076 407908 453082
rect 407856 453018 407908 453024
rect 407868 109041 407896 453018
rect 407854 109032 407910 109041
rect 407854 108967 407910 108976
rect 407762 17368 407818 17377
rect 407762 17303 407818 17312
rect 407960 17241 407988 454174
rect 408038 451616 408094 451625
rect 408038 451551 408094 451560
rect 408052 107506 408080 451551
rect 408314 450800 408370 450809
rect 408314 450735 408370 450744
rect 408130 450664 408186 450673
rect 408130 450599 408186 450608
rect 408144 107574 408172 450599
rect 408224 449608 408276 449614
rect 408224 449550 408276 449556
rect 408236 108905 408264 449550
rect 408328 109313 408356 450735
rect 408408 233912 408460 233918
rect 408408 233854 408460 233860
rect 408314 109304 408370 109313
rect 408314 109239 408370 109248
rect 408222 108896 408278 108905
rect 408222 108831 408278 108840
rect 408132 107568 408184 107574
rect 408132 107510 408184 107516
rect 408040 107500 408092 107506
rect 408040 107442 408092 107448
rect 407946 17232 408002 17241
rect 407946 17167 408002 17176
rect 407132 16546 407252 16574
rect 406384 3664 406436 3670
rect 406384 3606 406436 3612
rect 407224 480 407252 16546
rect 408420 3806 408448 233854
rect 409800 140078 409828 465122
rect 410524 454164 410576 454170
rect 410524 454106 410576 454112
rect 409880 247920 409932 247926
rect 409880 247862 409932 247868
rect 409788 140072 409840 140078
rect 409788 140014 409840 140020
rect 409892 16574 409920 247862
rect 410536 17814 410564 454106
rect 410708 453416 410760 453422
rect 410708 453358 410760 453364
rect 410614 451344 410670 451353
rect 410614 451279 410670 451288
rect 410628 106826 410656 451279
rect 410720 109070 410748 453358
rect 411076 450764 411128 450770
rect 411076 450706 411128 450712
rect 410984 450696 411036 450702
rect 410984 450638 411036 450644
rect 410892 450628 410944 450634
rect 410892 450570 410944 450576
rect 410800 450560 410852 450566
rect 410800 450502 410852 450508
rect 410708 109064 410760 109070
rect 410708 109006 410760 109012
rect 410812 108730 410840 450502
rect 410800 108724 410852 108730
rect 410800 108666 410852 108672
rect 410904 108594 410932 450570
rect 410892 108588 410944 108594
rect 410892 108530 410944 108536
rect 410996 108526 411024 450638
rect 410984 108520 411036 108526
rect 410984 108462 411036 108468
rect 411088 108458 411116 450706
rect 411180 141438 411208 466414
rect 411260 466404 411312 466410
rect 411260 466346 411312 466352
rect 411272 465118 411300 466346
rect 411260 465112 411312 465118
rect 411260 465054 411312 465060
rect 412548 465112 412600 465118
rect 412548 465054 412600 465060
rect 411904 244928 411956 244934
rect 411904 244870 411956 244876
rect 411168 141432 411220 141438
rect 411168 141374 411220 141380
rect 411076 108452 411128 108458
rect 411076 108394 411128 108400
rect 410616 106820 410668 106826
rect 410616 106762 410668 106768
rect 410524 17808 410576 17814
rect 410524 17750 410576 17756
rect 409892 16546 410840 16574
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 410812 480 410840 16546
rect 411916 4010 411944 244870
rect 412560 108662 412588 465054
rect 413376 453212 413428 453218
rect 413376 453154 413428 453160
rect 413284 451512 413336 451518
rect 413284 451454 413336 451460
rect 412548 108656 412600 108662
rect 412548 108598 412600 108604
rect 413296 108390 413324 451454
rect 413388 109342 413416 453154
rect 413468 450492 413520 450498
rect 413468 450434 413520 450440
rect 413376 109336 413428 109342
rect 413376 109278 413428 109284
rect 413480 108798 413508 450434
rect 413560 450424 413612 450430
rect 413560 450366 413612 450372
rect 413572 108866 413600 450366
rect 413652 450356 413704 450362
rect 413652 450298 413704 450304
rect 413664 109206 413692 450298
rect 413744 450288 413796 450294
rect 413744 450230 413796 450236
rect 413756 109274 413784 450230
rect 413940 144906 413968 469202
rect 414768 469198 414796 583442
rect 414860 471986 414888 584190
rect 415032 583432 415084 583438
rect 415032 583374 415084 583380
rect 414940 583296 414992 583302
rect 414940 583238 414992 583244
rect 414848 471980 414900 471986
rect 414848 471922 414900 471928
rect 414860 471442 414888 471922
rect 414848 471436 414900 471442
rect 414848 471378 414900 471384
rect 414756 469192 414808 469198
rect 414756 469134 414808 469140
rect 414768 468722 414796 469134
rect 414572 468716 414624 468722
rect 414572 468658 414624 468664
rect 414756 468716 414808 468722
rect 414756 468658 414808 468664
rect 414020 247852 414072 247858
rect 414020 247794 414072 247800
rect 413928 144900 413980 144906
rect 413928 144842 413980 144848
rect 413836 127628 413888 127634
rect 413836 127570 413888 127576
rect 413744 109268 413796 109274
rect 413744 109210 413796 109216
rect 413652 109200 413704 109206
rect 413652 109142 413704 109148
rect 413560 108860 413612 108866
rect 413560 108802 413612 108808
rect 413468 108792 413520 108798
rect 413468 108734 413520 108740
rect 413284 108384 413336 108390
rect 413284 108326 413336 108332
rect 411996 104644 412048 104650
rect 411996 104586 412048 104592
rect 412008 6254 412036 104586
rect 411996 6248 412048 6254
rect 411996 6190 412048 6196
rect 411904 4004 411956 4010
rect 411904 3946 411956 3952
rect 413848 3942 413876 127570
rect 414032 16574 414060 247794
rect 414584 113174 414612 468658
rect 414756 463004 414808 463010
rect 414756 462946 414808 462952
rect 414768 462466 414796 462946
rect 414756 462460 414808 462466
rect 414756 462402 414808 462408
rect 414664 124908 414716 124914
rect 414664 124850 414716 124856
rect 414492 113146 414612 113174
rect 414388 108248 414440 108254
rect 414388 108190 414440 108196
rect 414400 106026 414428 108190
rect 414492 106214 414520 113146
rect 414572 108044 414624 108050
rect 414572 107986 414624 107992
rect 414480 106208 414532 106214
rect 414480 106150 414532 106156
rect 414400 105998 414520 106026
rect 414584 106010 414612 107986
rect 414388 105596 414440 105602
rect 414388 105538 414440 105544
rect 414400 16998 414428 105538
rect 414492 17746 414520 105998
rect 414572 106004 414624 106010
rect 414572 105946 414624 105952
rect 414584 18494 414612 105946
rect 414572 18488 414624 18494
rect 414572 18430 414624 18436
rect 414480 17740 414532 17746
rect 414480 17682 414532 17688
rect 414388 16992 414440 16998
rect 414388 16934 414440 16940
rect 414032 16546 414336 16574
rect 413836 3936 413888 3942
rect 413836 3878 413888 3884
rect 414308 480 414336 16546
rect 414676 4146 414704 124850
rect 414768 106078 414796 462402
rect 414860 108254 414888 471378
rect 414952 466410 414980 583238
rect 415044 481642 415072 583374
rect 415872 535566 415900 586094
rect 415952 584656 416004 584662
rect 415952 584598 416004 584604
rect 415860 535560 415912 535566
rect 415860 535502 415912 535508
rect 415858 527232 415914 527241
rect 415858 527167 415914 527176
rect 415308 495236 415360 495242
rect 415308 495178 415360 495184
rect 415320 494902 415348 495178
rect 415308 494896 415360 494902
rect 415308 494838 415360 494844
rect 415216 490884 415268 490890
rect 415216 490826 415268 490832
rect 415228 490686 415256 490826
rect 415216 490680 415268 490686
rect 415216 490622 415268 490628
rect 415124 487212 415176 487218
rect 415124 487154 415176 487160
rect 415032 481636 415084 481642
rect 415032 481578 415084 481584
rect 415044 480282 415072 481578
rect 415032 480276 415084 480282
rect 415032 480218 415084 480224
rect 414940 466404 414992 466410
rect 414940 466346 414992 466352
rect 414848 108248 414900 108254
rect 414848 108190 414900 108196
rect 415044 106282 415072 480218
rect 415136 108186 415164 487154
rect 415124 108180 415176 108186
rect 415124 108122 415176 108128
rect 415228 108050 415256 490622
rect 415216 108044 415268 108050
rect 415216 107986 415268 107992
rect 415320 107930 415348 494838
rect 415872 465050 415900 527167
rect 415964 500206 415992 584598
rect 416056 500449 416084 586570
rect 416596 585064 416648 585070
rect 416596 585006 416648 585012
rect 416504 584996 416556 585002
rect 416504 584938 416556 584944
rect 416228 584928 416280 584934
rect 416228 584870 416280 584876
rect 416136 584588 416188 584594
rect 416136 584530 416188 584536
rect 416042 500440 416098 500449
rect 416042 500375 416098 500384
rect 415952 500200 416004 500206
rect 415952 500142 416004 500148
rect 416148 497418 416176 584530
rect 416240 500750 416268 584870
rect 416320 584792 416372 584798
rect 416320 584734 416372 584740
rect 416332 500886 416360 584734
rect 416412 584724 416464 584730
rect 416412 584666 416464 584672
rect 416424 500954 416452 584666
rect 416412 500948 416464 500954
rect 416412 500890 416464 500896
rect 416320 500880 416372 500886
rect 416320 500822 416372 500828
rect 416228 500744 416280 500750
rect 416228 500686 416280 500692
rect 416516 500682 416544 584938
rect 416504 500676 416556 500682
rect 416504 500618 416556 500624
rect 416608 500614 416636 585006
rect 416688 584860 416740 584866
rect 416688 584802 416740 584808
rect 416700 500818 416728 584802
rect 417160 536110 417188 625903
rect 417422 599992 417478 600001
rect 417422 599927 417478 599936
rect 417332 586288 417384 586294
rect 417332 586230 417384 586236
rect 417240 583364 417292 583370
rect 417240 583306 417292 583312
rect 417148 536104 417200 536110
rect 417148 536046 417200 536052
rect 417160 535945 417188 536046
rect 417146 535936 417202 535945
rect 417146 535871 417202 535880
rect 416780 535560 416832 535566
rect 416780 535502 416832 535508
rect 416688 500812 416740 500818
rect 416688 500754 416740 500760
rect 416596 500608 416648 500614
rect 416596 500550 416648 500556
rect 416136 497412 416188 497418
rect 416136 497354 416188 497360
rect 416686 494048 416742 494057
rect 416686 493983 416742 493992
rect 416700 492726 416728 493983
rect 416688 492720 416740 492726
rect 416688 492662 416740 492668
rect 415860 465044 415912 465050
rect 415860 464986 415912 464992
rect 416044 451716 416096 451722
rect 416044 451658 416096 451664
rect 415400 246356 415452 246362
rect 415400 246298 415452 246304
rect 415412 117978 415440 246298
rect 415952 123480 416004 123486
rect 415952 123422 416004 123428
rect 415400 117972 415452 117978
rect 415400 117914 415452 117920
rect 415136 107902 415348 107930
rect 415136 107030 415164 107902
rect 415124 107024 415176 107030
rect 415124 106966 415176 106972
rect 415032 106276 415084 106282
rect 415032 106218 415084 106224
rect 414756 106072 414808 106078
rect 414756 106014 414808 106020
rect 414768 105602 414796 106014
rect 414756 105596 414808 105602
rect 414756 105538 414808 105544
rect 414940 104576 414992 104582
rect 414940 104518 414992 104524
rect 414756 104508 414808 104514
rect 414756 104450 414808 104456
rect 414664 4140 414716 4146
rect 414664 4082 414716 4088
rect 414768 3505 414796 104450
rect 414848 104440 414900 104446
rect 414848 104382 414900 104388
rect 414754 3496 414810 3505
rect 414754 3431 414810 3440
rect 414860 3398 414888 104382
rect 414848 3392 414900 3398
rect 414952 3369 414980 104518
rect 415136 18426 415164 106966
rect 415308 106208 415360 106214
rect 415308 106150 415360 106156
rect 415320 19310 415348 106150
rect 415308 19304 415360 19310
rect 415308 19246 415360 19252
rect 415124 18420 415176 18426
rect 415124 18362 415176 18368
rect 414848 3334 414900 3340
rect 414938 3360 414994 3369
rect 414938 3295 414994 3304
rect 415964 3194 415992 123422
rect 416056 18970 416084 451658
rect 416320 450900 416372 450906
rect 416320 450842 416372 450848
rect 416136 450152 416188 450158
rect 416136 450094 416188 450100
rect 416148 109614 416176 450094
rect 416228 450016 416280 450022
rect 416228 449958 416280 449964
rect 416136 109608 416188 109614
rect 416136 109550 416188 109556
rect 416240 109478 416268 449958
rect 416228 109472 416280 109478
rect 416228 109414 416280 109420
rect 416332 109410 416360 450842
rect 416412 450084 416464 450090
rect 416412 450026 416464 450032
rect 416424 109546 416452 450026
rect 416504 180124 416556 180130
rect 416504 180066 416556 180072
rect 416412 109540 416464 109546
rect 416412 109482 416464 109488
rect 416320 109404 416372 109410
rect 416320 109346 416372 109352
rect 416136 108656 416188 108662
rect 416136 108598 416188 108604
rect 416148 107778 416176 108598
rect 416412 108180 416464 108186
rect 416412 108122 416464 108128
rect 416424 107846 416452 108122
rect 416412 107840 416464 107846
rect 416412 107782 416464 107788
rect 416136 107772 416188 107778
rect 416136 107714 416188 107720
rect 416044 18964 416096 18970
rect 416044 18906 416096 18912
rect 416148 16590 416176 107714
rect 416320 107704 416372 107710
rect 416320 107646 416372 107652
rect 416228 106276 416280 106282
rect 416228 106218 416280 106224
rect 416240 105602 416268 106218
rect 416228 105596 416280 105602
rect 416228 105538 416280 105544
rect 416240 19242 416268 105538
rect 416332 19786 416360 107646
rect 416320 19780 416372 19786
rect 416320 19722 416372 19728
rect 416228 19236 416280 19242
rect 416228 19178 416280 19184
rect 416424 19174 416452 107782
rect 416412 19168 416464 19174
rect 416412 19110 416464 19116
rect 416136 16584 416188 16590
rect 416136 16526 416188 16532
rect 416516 3534 416544 180066
rect 416596 126268 416648 126274
rect 416596 126210 416648 126216
rect 416608 4078 416636 126210
rect 416700 107522 416728 492662
rect 416792 492658 416820 535502
rect 416870 531040 416926 531049
rect 416870 530975 416926 530984
rect 416884 530670 416912 530975
rect 416872 530664 416924 530670
rect 416872 530606 416924 530612
rect 416964 530596 417016 530602
rect 416964 530538 417016 530544
rect 416976 529961 417004 530538
rect 416962 529952 417018 529961
rect 416962 529887 417018 529896
rect 416870 509960 416926 509969
rect 416870 509895 416872 509904
rect 416924 509895 416926 509904
rect 416872 509866 416924 509872
rect 417252 496874 417280 583306
rect 417344 496942 417372 586230
rect 417436 509969 417464 599927
rect 417528 537538 417556 626855
rect 418066 623792 418122 623801
rect 418066 623727 418122 623736
rect 417974 621072 418030 621081
rect 417974 621007 418030 621016
rect 417606 619984 417662 619993
rect 417606 619919 417662 619928
rect 417516 537532 417568 537538
rect 417516 537474 417568 537480
rect 417528 536897 417556 537474
rect 417514 536888 417570 536897
rect 417514 536823 417570 536832
rect 417514 533760 417570 533769
rect 417514 533695 417516 533704
rect 417568 533695 417570 533704
rect 417516 533666 417568 533672
rect 417620 530602 417648 619919
rect 417792 591388 417844 591394
rect 417792 591330 417844 591336
rect 417700 587172 417752 587178
rect 417700 587114 417752 587120
rect 417712 586945 417740 587114
rect 417698 586936 417754 586945
rect 417698 586871 417754 586880
rect 417804 586498 417832 591330
rect 417792 586492 417844 586498
rect 417792 586434 417844 586440
rect 417700 586424 417752 586430
rect 417700 586366 417752 586372
rect 417608 530596 417660 530602
rect 417608 530538 417660 530544
rect 417422 509960 417478 509969
rect 417422 509895 417478 509904
rect 417422 508056 417478 508065
rect 417422 507991 417478 508000
rect 417332 496936 417384 496942
rect 417332 496878 417384 496884
rect 417240 496868 417292 496874
rect 417240 496810 417292 496816
rect 416780 492652 416832 492658
rect 416780 492594 416832 492600
rect 417436 474230 417464 507991
rect 417424 474224 417476 474230
rect 417424 474166 417476 474172
rect 417712 470558 417740 586366
rect 417804 508337 417832 586434
rect 417884 535492 417936 535498
rect 417884 535434 417936 535440
rect 417790 508328 417846 508337
rect 417790 508263 417846 508272
rect 417804 507890 417832 508263
rect 417792 507884 417844 507890
rect 417792 507826 417844 507832
rect 417792 492652 417844 492658
rect 417792 492594 417844 492600
rect 417804 491366 417832 492594
rect 417792 491360 417844 491366
rect 417792 491302 417844 491308
rect 417700 470552 417752 470558
rect 417700 470494 417752 470500
rect 417712 469334 417740 470494
rect 417700 469328 417752 469334
rect 417700 469270 417752 469276
rect 417424 465044 417476 465050
rect 417424 464986 417476 464992
rect 417436 464506 417464 464986
rect 417424 464500 417476 464506
rect 417424 464442 417476 464448
rect 417436 463729 417464 464442
rect 417422 463720 417478 463729
rect 417422 463655 417478 463664
rect 417424 452328 417476 452334
rect 417424 452270 417476 452276
rect 416778 146976 416834 146985
rect 416778 146911 416780 146920
rect 416832 146911 416834 146920
rect 417330 146976 417386 146985
rect 417330 146911 417386 146920
rect 416780 146882 416832 146888
rect 417148 144900 417200 144906
rect 417148 144842 417200 144848
rect 417160 143857 417188 144842
rect 417146 143848 417202 143857
rect 417146 143783 417202 143792
rect 416780 141432 416832 141438
rect 416780 141374 416832 141380
rect 416792 141137 416820 141374
rect 416778 141128 416834 141137
rect 416778 141063 416834 141072
rect 416780 140072 416832 140078
rect 416778 140040 416780 140049
rect 416832 140040 416834 140049
rect 416778 139975 416834 139984
rect 417160 137358 417188 143783
rect 417238 140040 417294 140049
rect 417238 139975 417294 139984
rect 417148 137352 417200 137358
rect 417148 137294 417200 137300
rect 417146 120048 417202 120057
rect 417146 119983 417202 119992
rect 416700 107494 417096 107522
rect 417068 106418 417096 107494
rect 417056 106412 417108 106418
rect 417056 106354 417108 106360
rect 416780 28960 416832 28966
rect 416780 28902 416832 28908
rect 416792 28121 416820 28902
rect 416870 28384 416926 28393
rect 416870 28319 416926 28328
rect 416884 28286 416912 28319
rect 416872 28280 416924 28286
rect 416872 28222 416924 28228
rect 416778 28112 416834 28121
rect 416778 28047 416834 28056
rect 417068 17474 417096 106354
rect 417160 104854 417188 119983
rect 417148 104848 417200 104854
rect 417148 104790 417200 104796
rect 417252 50017 417280 139975
rect 417344 56953 417372 146911
rect 417436 118153 417464 452270
rect 417514 141128 417570 141137
rect 417514 141063 417570 141072
rect 417422 118144 417478 118153
rect 417422 118079 417478 118088
rect 417424 104848 417476 104854
rect 417424 104790 417476 104796
rect 417330 56944 417386 56953
rect 417330 56879 417386 56888
rect 417238 50008 417294 50017
rect 417238 49943 417294 49952
rect 417436 30025 417464 104790
rect 417528 51105 417556 141063
rect 417608 137352 417660 137358
rect 417608 137294 417660 137300
rect 417620 53825 417648 137294
rect 417712 106214 417740 469270
rect 417804 120222 417832 491302
rect 417896 488510 417924 535434
rect 417988 531049 418016 621007
rect 418080 533769 418108 623727
rect 419446 598362 419502 598371
rect 419446 598297 419502 598306
rect 419460 591394 419488 598297
rect 419448 591388 419500 591394
rect 419448 591330 419500 591336
rect 436282 587888 436338 587897
rect 436282 587823 436338 587832
rect 438122 587888 438178 587897
rect 438122 587823 438178 587832
rect 439594 587888 439650 587897
rect 439594 587823 439650 587832
rect 441618 587888 441674 587897
rect 441618 587823 441674 587832
rect 443090 587888 443146 587897
rect 443090 587823 443146 587832
rect 444194 587888 444250 587897
rect 444194 587823 444250 587832
rect 445666 587888 445722 587897
rect 445666 587823 445722 587832
rect 446494 587888 446550 587897
rect 446494 587823 446550 587832
rect 447322 587888 447378 587897
rect 447322 587823 447378 587832
rect 448518 587888 448574 587897
rect 448518 587823 448574 587832
rect 449898 587888 449954 587897
rect 449898 587823 449954 587832
rect 450634 587888 450690 587897
rect 450634 587823 450690 587832
rect 453578 587888 453634 587897
rect 453578 587823 453634 587832
rect 454590 587888 454646 587897
rect 454590 587823 454646 587832
rect 456062 587888 456118 587897
rect 456062 587823 456118 587832
rect 456798 587888 456854 587897
rect 456798 587823 456854 587832
rect 457258 587888 457314 587897
rect 457258 587823 457314 587832
rect 471242 587888 471298 587897
rect 471242 587823 471298 587832
rect 472162 587888 472218 587897
rect 473358 587888 473414 587897
rect 472162 587823 472218 587832
rect 473268 587852 473320 587858
rect 419170 587616 419226 587625
rect 419170 587551 419226 587560
rect 418710 587480 418766 587489
rect 418710 587415 418766 587424
rect 418620 586220 418672 586226
rect 418620 586162 418672 586168
rect 418632 535498 418660 586162
rect 418620 535492 418672 535498
rect 418620 535434 418672 535440
rect 418066 533760 418122 533769
rect 418066 533695 418122 533704
rect 417974 531040 418030 531049
rect 417974 530975 418030 530984
rect 418724 500274 418752 587415
rect 418986 587344 419042 587353
rect 418986 587279 419042 587288
rect 418804 586968 418856 586974
rect 418804 586910 418856 586916
rect 418712 500268 418764 500274
rect 418712 500210 418764 500216
rect 417976 497548 418028 497554
rect 417976 497490 418028 497496
rect 417988 496874 418016 497490
rect 418068 497480 418120 497486
rect 418068 497422 418120 497428
rect 418080 496942 418108 497422
rect 418068 496936 418120 496942
rect 418068 496878 418120 496884
rect 417976 496868 418028 496874
rect 417976 496810 418028 496816
rect 417884 488504 417936 488510
rect 417884 488446 417936 488452
rect 417896 487218 417924 488446
rect 417884 487212 417936 487218
rect 417884 487154 417936 487160
rect 417884 484356 417936 484362
rect 417884 484298 417936 484304
rect 417896 483886 417924 484298
rect 417884 483880 417936 483886
rect 417884 483822 417936 483828
rect 417792 120216 417844 120222
rect 417792 120158 417844 120164
rect 417790 118416 417846 118425
rect 417790 118351 417846 118360
rect 417804 117978 417832 118351
rect 417792 117972 417844 117978
rect 417792 117914 417844 117920
rect 417804 106282 417832 117914
rect 417896 107438 417924 483822
rect 417988 109750 418016 496810
rect 417976 109744 418028 109750
rect 417976 109686 418028 109692
rect 417884 107432 417936 107438
rect 417884 107374 417936 107380
rect 417792 106276 417844 106282
rect 417792 106218 417844 106224
rect 417700 106208 417752 106214
rect 417700 106150 417752 106156
rect 417606 53816 417662 53825
rect 417606 53751 417662 53760
rect 417514 51096 417570 51105
rect 417514 51031 417570 51040
rect 417422 30016 417478 30025
rect 417422 29951 417478 29960
rect 417804 28393 417832 106218
rect 417790 28384 417846 28393
rect 417790 28319 417846 28328
rect 417056 17468 417108 17474
rect 417056 17410 417108 17416
rect 417988 16386 418016 109686
rect 418080 107982 418108 496878
rect 418710 496768 418766 496777
rect 418710 496703 418766 496712
rect 418160 495576 418212 495582
rect 418160 495518 418212 495524
rect 418068 107976 418120 107982
rect 418068 107918 418120 107924
rect 418172 107710 418200 495518
rect 418724 495514 418752 496703
rect 418712 495508 418764 495514
rect 418712 495450 418764 495456
rect 418528 111104 418580 111110
rect 418528 111046 418580 111052
rect 418436 107976 418488 107982
rect 418436 107918 418488 107924
rect 418344 107908 418396 107914
rect 418344 107850 418396 107856
rect 418160 107704 418212 107710
rect 418160 107646 418212 107652
rect 418066 107536 418122 107545
rect 418066 107471 418122 107480
rect 418080 106486 418108 107471
rect 418068 106480 418120 106486
rect 418068 106422 418120 106428
rect 418080 17406 418108 106422
rect 418068 17400 418120 17406
rect 418068 17342 418120 17348
rect 418356 16522 418384 107850
rect 418448 22438 418476 107918
rect 418436 22432 418488 22438
rect 418436 22374 418488 22380
rect 418434 19136 418490 19145
rect 418434 19071 418490 19080
rect 418448 16930 418476 19071
rect 418436 16924 418488 16930
rect 418436 16866 418488 16872
rect 418344 16516 418396 16522
rect 418344 16458 418396 16464
rect 417976 16380 418028 16386
rect 417976 16322 418028 16328
rect 416596 4072 416648 4078
rect 416596 4014 416648 4020
rect 416504 3528 416556 3534
rect 416504 3470 416556 3476
rect 417884 3528 417936 3534
rect 417884 3470 417936 3476
rect 415952 3188 416004 3194
rect 415952 3130 416004 3136
rect 417896 480 417924 3470
rect 418540 3262 418568 111046
rect 418724 107234 418752 495450
rect 418816 468654 418844 586910
rect 418896 585132 418948 585138
rect 418896 585074 418948 585080
rect 418908 500546 418936 585074
rect 418896 500540 418948 500546
rect 418896 500482 418948 500488
rect 419000 500342 419028 587279
rect 419080 584316 419132 584322
rect 419080 584258 419132 584264
rect 419092 500410 419120 584258
rect 419184 500585 419212 587551
rect 420000 587512 420052 587518
rect 420000 587454 420052 587460
rect 419908 587308 419960 587314
rect 419908 587250 419960 587256
rect 419816 587240 419868 587246
rect 419816 587182 419868 587188
rect 419724 586696 419776 586702
rect 419724 586638 419776 586644
rect 419356 586356 419408 586362
rect 419356 586298 419408 586304
rect 419264 584384 419316 584390
rect 419264 584326 419316 584332
rect 419170 500576 419226 500585
rect 419170 500511 419226 500520
rect 419276 500478 419304 584326
rect 419264 500472 419316 500478
rect 419264 500414 419316 500420
rect 419080 500404 419132 500410
rect 419080 500346 419132 500352
rect 418988 500336 419040 500342
rect 418988 500278 419040 500284
rect 419368 480214 419396 586298
rect 419448 583568 419500 583574
rect 419448 583510 419500 583516
rect 419460 496738 419488 583510
rect 419736 498846 419764 586638
rect 419724 498840 419776 498846
rect 419724 498782 419776 498788
rect 419828 497622 419856 587182
rect 419920 497690 419948 587250
rect 419908 497684 419960 497690
rect 419908 497626 419960 497632
rect 419816 497616 419868 497622
rect 419816 497558 419868 497564
rect 420012 496806 420040 587454
rect 436296 584905 436324 587823
rect 438136 587314 438164 587823
rect 438124 587308 438176 587314
rect 438124 587250 438176 587256
rect 439608 587246 439636 587823
rect 439596 587240 439648 587246
rect 439596 587182 439648 587188
rect 441632 587178 441660 587823
rect 441620 587172 441672 587178
rect 441620 587114 441672 587120
rect 443104 587110 443132 587823
rect 443092 587104 443144 587110
rect 443092 587046 443144 587052
rect 444208 587042 444236 587823
rect 445680 587314 445708 587823
rect 445668 587308 445720 587314
rect 445668 587250 445720 587256
rect 444196 587036 444248 587042
rect 444196 586978 444248 586984
rect 445680 586906 445708 587250
rect 445668 586900 445720 586906
rect 445668 586842 445720 586848
rect 446508 586838 446536 587823
rect 447336 586906 447364 587823
rect 448532 587110 448560 587823
rect 449912 587178 449940 587823
rect 449900 587172 449952 587178
rect 449900 587114 449952 587120
rect 448520 587104 448572 587110
rect 448520 587046 448572 587052
rect 447324 586900 447376 586906
rect 447324 586842 447376 586848
rect 445760 586832 445812 586838
rect 445760 586774 445812 586780
rect 446496 586832 446548 586838
rect 446496 586774 446548 586780
rect 436282 584896 436338 584905
rect 436282 584831 436338 584840
rect 445772 583574 445800 586774
rect 445760 583568 445812 583574
rect 445760 583510 445812 583516
rect 447336 583506 447364 586842
rect 447324 583500 447376 583506
rect 447324 583442 447376 583448
rect 448532 583438 448560 587046
rect 449912 586430 449940 587114
rect 450648 587042 450676 587823
rect 452382 587752 452438 587761
rect 452382 587687 452438 587696
rect 453486 587752 453542 587761
rect 453486 587687 453542 587696
rect 450820 587172 450872 587178
rect 450820 587114 450872 587120
rect 450636 587036 450688 587042
rect 450636 586978 450688 586984
rect 450832 586974 450860 587114
rect 450820 586968 450872 586974
rect 450820 586910 450872 586916
rect 451370 586936 451426 586945
rect 451370 586871 451426 586880
rect 451384 586838 451412 586871
rect 451372 586832 451424 586838
rect 451372 586774 451424 586780
rect 451280 586764 451332 586770
rect 451280 586706 451332 586712
rect 449900 586424 449952 586430
rect 449900 586366 449952 586372
rect 451292 586294 451320 586706
rect 451280 586288 451332 586294
rect 451280 586230 451332 586236
rect 448520 583432 448572 583438
rect 448520 583374 448572 583380
rect 451384 583370 451412 586774
rect 452396 586770 452424 587687
rect 452660 587376 452712 587382
rect 452660 587318 452712 587324
rect 452384 586764 452436 586770
rect 452384 586706 452436 586712
rect 452672 586702 452700 587318
rect 453500 586702 453528 587687
rect 452660 586696 452712 586702
rect 452660 586638 452712 586644
rect 452752 586696 452804 586702
rect 452752 586638 452804 586644
rect 453488 586696 453540 586702
rect 453488 586638 453540 586644
rect 452764 586362 452792 586638
rect 453592 586634 453620 587823
rect 454604 587382 454632 587823
rect 456076 587586 456104 587823
rect 456154 587752 456210 587761
rect 456154 587687 456210 587696
rect 456064 587580 456116 587586
rect 456064 587522 456116 587528
rect 454592 587376 454644 587382
rect 454592 587318 454644 587324
rect 456168 586702 456196 587687
rect 456812 586945 456840 587823
rect 456798 586936 456854 586945
rect 456798 586871 456854 586880
rect 456156 586696 456208 586702
rect 456156 586638 456208 586644
rect 453580 586628 453632 586634
rect 453580 586570 453632 586576
rect 452752 586356 452804 586362
rect 452752 586298 452804 586304
rect 456168 586226 456196 586638
rect 456156 586220 456208 586226
rect 456156 586162 456208 586168
rect 456812 586158 456840 586871
rect 456800 586152 456852 586158
rect 456800 586094 456852 586100
rect 457272 584254 457300 587823
rect 458270 587752 458326 587761
rect 458270 587687 458326 587696
rect 460662 587752 460718 587761
rect 460662 587687 460718 587696
rect 460938 587752 460994 587761
rect 460938 587687 460994 587696
rect 461582 587752 461638 587761
rect 461582 587687 461638 587696
rect 462318 587752 462374 587761
rect 462318 587687 462374 587696
rect 463882 587752 463938 587761
rect 463882 587687 463938 587696
rect 465078 587752 465134 587761
rect 465078 587687 465134 587696
rect 466274 587752 466330 587761
rect 466274 587687 466330 587696
rect 467562 587752 467618 587761
rect 467562 587687 467618 587696
rect 468666 587752 468722 587761
rect 468666 587687 468722 587696
rect 469770 587752 469826 587761
rect 469770 587687 469826 587696
rect 458178 587208 458234 587217
rect 458178 587143 458234 587152
rect 458192 586566 458220 587143
rect 458284 586566 458312 587687
rect 459744 587512 459796 587518
rect 459744 587454 459796 587460
rect 459756 587178 459784 587454
rect 460676 587178 460704 587687
rect 459744 587172 459796 587178
rect 459744 587114 459796 587120
rect 460664 587172 460716 587178
rect 460664 587114 460716 587120
rect 458180 586560 458232 586566
rect 458180 586502 458232 586508
rect 458272 586560 458324 586566
rect 458272 586502 458324 586508
rect 457260 584248 457312 584254
rect 457260 584190 457312 584196
rect 458284 583370 458312 586502
rect 460952 584769 460980 587687
rect 461596 587450 461624 587687
rect 461584 587444 461636 587450
rect 461584 587386 461636 587392
rect 462332 586090 462360 587687
rect 463896 587314 463924 587687
rect 463884 587308 463936 587314
rect 463884 587250 463936 587256
rect 462780 587240 462832 587246
rect 462778 587208 462780 587217
rect 462832 587208 462834 587217
rect 462778 587143 462834 587152
rect 462320 586084 462372 586090
rect 462320 586026 462372 586032
rect 460938 584760 460994 584769
rect 460938 584695 460994 584704
rect 465092 584633 465120 587687
rect 465170 587208 465226 587217
rect 465170 587143 465226 587152
rect 465184 586906 465212 587143
rect 466288 587042 466316 587687
rect 467576 587110 467604 587687
rect 467564 587104 467616 587110
rect 467564 587046 467616 587052
rect 466276 587036 466328 587042
rect 466276 586978 466328 586984
rect 468680 586974 468708 587687
rect 468668 586968 468720 586974
rect 468668 586910 468720 586916
rect 465172 586900 465224 586906
rect 465172 586842 465224 586848
rect 469784 586838 469812 587687
rect 469772 586832 469824 586838
rect 469772 586774 469824 586780
rect 471256 586770 471284 587823
rect 471244 586764 471296 586770
rect 471244 586706 471296 586712
rect 472176 586634 472204 587823
rect 473358 587823 473414 587832
rect 473634 587888 473690 587897
rect 473634 587823 473690 587832
rect 476946 587888 477002 587897
rect 476946 587823 476948 587832
rect 473268 587794 473320 587800
rect 473280 587761 473308 587794
rect 473266 587752 473322 587761
rect 473266 587687 473322 587696
rect 473372 587382 473400 587823
rect 473360 587376 473412 587382
rect 473360 587318 473412 587324
rect 473648 586702 473676 587823
rect 477000 587823 477002 587832
rect 478050 587888 478106 587897
rect 478050 587823 478106 587832
rect 479154 587888 479210 587897
rect 479154 587823 479210 587832
rect 480258 587888 480314 587897
rect 480258 587823 480314 587832
rect 483018 587888 483074 587897
rect 483018 587823 483074 587832
rect 485778 587888 485834 587897
rect 485778 587823 485834 587832
rect 487158 587888 487214 587897
rect 487158 587823 487214 587832
rect 492678 587888 492734 587897
rect 492678 587823 492734 587832
rect 495438 587888 495494 587897
rect 495438 587823 495494 587832
rect 498198 587888 498254 587897
rect 498198 587823 498254 587832
rect 500958 587888 501014 587897
rect 500958 587823 501014 587832
rect 502338 587888 502394 587897
rect 502338 587823 502394 587832
rect 505098 587888 505154 587897
rect 505098 587823 505154 587832
rect 507858 587888 507914 587897
rect 507858 587823 507914 587832
rect 510618 587888 510674 587897
rect 510618 587823 510674 587832
rect 513378 587888 513434 587897
rect 513378 587823 513434 587832
rect 514758 587888 514814 587897
rect 514758 587823 514814 587832
rect 520278 587888 520334 587897
rect 523314 587888 523370 587897
rect 520278 587823 520334 587832
rect 522396 587852 522448 587858
rect 476948 587794 477000 587800
rect 473636 586696 473688 586702
rect 473636 586638 473688 586644
rect 472164 586628 472216 586634
rect 472164 586570 472216 586576
rect 474096 586628 474148 586634
rect 474096 586570 474148 586576
rect 470598 586528 470654 586537
rect 470598 586463 470654 586472
rect 470612 586022 470640 586463
rect 470600 586016 470652 586022
rect 470600 585958 470652 585964
rect 465078 584624 465134 584633
rect 465078 584559 465134 584568
rect 474108 584526 474136 586570
rect 478064 586566 478092 587823
rect 479168 587178 479196 587823
rect 479156 587172 479208 587178
rect 479156 587114 479208 587120
rect 478052 586560 478104 586566
rect 478052 586502 478104 586508
rect 474096 584520 474148 584526
rect 474096 584462 474148 584468
rect 480272 584322 480300 587823
rect 483032 584390 483060 587823
rect 485792 585138 485820 587823
rect 485780 585132 485832 585138
rect 485780 585074 485832 585080
rect 487172 585070 487200 587823
rect 489918 586528 489974 586537
rect 489918 586463 489974 586472
rect 487160 585064 487212 585070
rect 487160 585006 487212 585012
rect 489932 585002 489960 586463
rect 489920 584996 489972 585002
rect 489920 584938 489972 584944
rect 492692 584934 492720 587823
rect 492680 584928 492732 584934
rect 492680 584870 492732 584876
rect 495452 584866 495480 587823
rect 495440 584860 495492 584866
rect 495440 584802 495492 584808
rect 498212 584798 498240 587823
rect 498200 584792 498252 584798
rect 498200 584734 498252 584740
rect 500972 584730 501000 587823
rect 500960 584724 501012 584730
rect 500960 584666 501012 584672
rect 502352 584662 502380 587823
rect 502340 584656 502392 584662
rect 502340 584598 502392 584604
rect 505112 584594 505140 587823
rect 505100 584588 505152 584594
rect 505100 584530 505152 584536
rect 507872 584497 507900 587823
rect 507858 584488 507914 584497
rect 510632 584458 510660 587823
rect 513392 585954 513420 587823
rect 513380 585948 513432 585954
rect 513380 585890 513432 585896
rect 507858 584423 507914 584432
rect 510620 584452 510672 584458
rect 510620 584394 510672 584400
rect 483020 584384 483072 584390
rect 514772 584361 514800 587823
rect 520292 585818 520320 587823
rect 523314 587823 523370 587832
rect 525890 587888 525946 587897
rect 525890 587823 525892 587832
rect 522396 587794 522448 587800
rect 522408 585886 522436 587794
rect 523328 586634 523356 587823
rect 525944 587823 525946 587832
rect 525892 587794 525944 587800
rect 523316 586628 523368 586634
rect 523316 586570 523368 586576
rect 557552 586498 557580 674834
rect 565084 670744 565136 670750
rect 580172 670744 580224 670750
rect 565084 670686 565136 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 558918 668672 558974 668681
rect 558918 668607 558974 668616
rect 558184 590708 558236 590714
rect 558184 590650 558236 590656
rect 550824 586492 550876 586498
rect 550824 586434 550876 586440
rect 557540 586492 557592 586498
rect 557540 586434 557592 586440
rect 522396 585880 522448 585886
rect 522396 585822 522448 585828
rect 520280 585812 520332 585818
rect 520280 585754 520332 585760
rect 550836 585313 550864 586434
rect 550822 585304 550878 585313
rect 550822 585239 550878 585248
rect 483020 584326 483072 584332
rect 514758 584352 514814 584361
rect 480260 584316 480312 584322
rect 514758 584287 514814 584296
rect 480260 584258 480312 584264
rect 451372 583364 451424 583370
rect 451372 583306 451424 583312
rect 458272 583364 458324 583370
rect 458272 583306 458324 583312
rect 558196 498914 558224 590650
rect 558932 579193 558960 668607
rect 563704 616888 563756 616894
rect 563704 616830 563756 616836
rect 558918 579184 558974 579193
rect 558918 579119 558974 579128
rect 558276 510672 558328 510678
rect 558276 510614 558328 510620
rect 558184 498908 558236 498914
rect 558184 498850 558236 498856
rect 454592 498840 454644 498846
rect 454592 498782 454644 498788
rect 454604 498166 454632 498782
rect 454592 498160 454644 498166
rect 441618 498128 441674 498137
rect 441618 498063 441674 498072
rect 445298 498128 445354 498137
rect 445298 498063 445354 498072
rect 449162 498128 449218 498137
rect 449162 498063 449218 498072
rect 451278 498128 451334 498137
rect 451278 498063 451334 498072
rect 452382 498128 452438 498137
rect 452382 498063 452438 498072
rect 454590 498128 454592 498137
rect 473360 498160 473412 498166
rect 454644 498128 454646 498137
rect 454590 498063 454646 498072
rect 455510 498128 455566 498137
rect 455510 498063 455566 498072
rect 469218 498128 469274 498137
rect 469218 498063 469274 498072
rect 473358 498128 473360 498137
rect 473412 498128 473414 498137
rect 473358 498063 473414 498072
rect 473542 498128 473598 498137
rect 473542 498063 473598 498072
rect 480534 498128 480590 498137
rect 480534 498063 480590 498072
rect 494702 498128 494758 498137
rect 494702 498063 494758 498072
rect 504362 498128 504418 498137
rect 504362 498063 504418 498072
rect 512642 498128 512698 498137
rect 512642 498063 512698 498072
rect 519542 498128 519598 498137
rect 519542 498063 519598 498072
rect 436190 497992 436246 498001
rect 436190 497927 436246 497936
rect 436204 497049 436232 497927
rect 437480 497684 437532 497690
rect 437480 497626 437532 497632
rect 436190 497040 436246 497049
rect 436190 496975 436246 496984
rect 436098 496904 436154 496913
rect 420736 496868 420788 496874
rect 436098 496839 436100 496848
rect 420736 496810 420788 496816
rect 436152 496839 436154 496848
rect 436100 496810 436152 496816
rect 420000 496800 420052 496806
rect 420748 496777 420776 496810
rect 420000 496742 420052 496748
rect 420734 496768 420790 496777
rect 419448 496732 419500 496738
rect 419448 496674 419500 496680
rect 420012 495582 420040 496742
rect 420734 496703 420790 496712
rect 420000 495576 420052 495582
rect 420000 495518 420052 495524
rect 419356 480208 419408 480214
rect 419356 480150 419408 480156
rect 419368 479534 419396 480150
rect 419356 479528 419408 479534
rect 419356 479470 419408 479476
rect 420000 479528 420052 479534
rect 420000 479470 420052 479476
rect 418804 468648 418856 468654
rect 418804 468590 418856 468596
rect 419448 463140 419500 463146
rect 419448 463082 419500 463088
rect 419460 462398 419488 463082
rect 419448 462392 419500 462398
rect 419448 462334 419500 462340
rect 418804 453008 418856 453014
rect 418804 452950 418856 452956
rect 418816 107273 418844 452950
rect 418896 452396 418948 452402
rect 418896 452338 418948 452344
rect 418908 108662 418936 452338
rect 419460 451274 419488 462334
rect 419632 456340 419684 456346
rect 419632 456282 419684 456288
rect 419540 456272 419592 456278
rect 419540 456214 419592 456220
rect 419552 455938 419580 456214
rect 419644 456142 419672 456282
rect 419724 456204 419776 456210
rect 419724 456146 419776 456152
rect 419632 456136 419684 456142
rect 419632 456078 419684 456084
rect 419540 455932 419592 455938
rect 419540 455874 419592 455880
rect 419368 451246 419488 451274
rect 418988 450220 419040 450226
rect 418988 450162 419040 450168
rect 419000 109682 419028 450162
rect 419264 120216 419316 120222
rect 419264 120158 419316 120164
rect 419080 112464 419132 112470
rect 419080 112406 419132 112412
rect 418988 109676 419040 109682
rect 418988 109618 419040 109624
rect 418896 108656 418948 108662
rect 418896 108598 418948 108604
rect 418896 107704 418948 107710
rect 418896 107646 418948 107652
rect 418908 107370 418936 107646
rect 418896 107364 418948 107370
rect 418896 107306 418948 107312
rect 418802 107264 418858 107273
rect 418712 107228 418764 107234
rect 418802 107199 418858 107208
rect 418712 107170 418764 107176
rect 418620 106208 418672 106214
rect 418620 106150 418672 106156
rect 418632 105670 418660 106150
rect 418620 105664 418672 105670
rect 418620 105606 418672 105612
rect 418632 22522 418660 105606
rect 418724 22642 418752 107170
rect 418896 106956 418948 106962
rect 418896 106898 418948 106904
rect 418804 104168 418856 104174
rect 418804 104110 418856 104116
rect 418712 22636 418764 22642
rect 418712 22578 418764 22584
rect 418632 22494 418752 22522
rect 418620 22432 418672 22438
rect 418620 22374 418672 22380
rect 418632 16250 418660 22374
rect 418724 18562 418752 22494
rect 418712 18556 418764 18562
rect 418712 18498 418764 18504
rect 418620 16244 418672 16250
rect 418620 16186 418672 16192
rect 418816 3874 418844 104110
rect 418804 3868 418856 3874
rect 418804 3810 418856 3816
rect 418908 3738 418936 106898
rect 418988 106888 419040 106894
rect 418988 106830 419040 106836
rect 419000 17134 419028 106830
rect 418988 17128 419040 17134
rect 418988 17070 419040 17076
rect 418896 3732 418948 3738
rect 418896 3674 418948 3680
rect 419092 3330 419120 112406
rect 419276 107914 419304 120158
rect 419264 107908 419316 107914
rect 419264 107850 419316 107856
rect 419264 107432 419316 107438
rect 419264 107374 419316 107380
rect 419276 106350 419304 107374
rect 419368 106894 419396 451246
rect 419736 107098 419764 456146
rect 419908 456136 419960 456142
rect 419908 456078 419960 456084
rect 419816 455932 419868 455938
rect 419816 455874 419868 455880
rect 419828 107166 419856 455874
rect 419816 107160 419868 107166
rect 419816 107102 419868 107108
rect 419724 107092 419776 107098
rect 419724 107034 419776 107040
rect 419356 106888 419408 106894
rect 419356 106830 419408 106836
rect 419264 106344 419316 106350
rect 419264 106286 419316 106292
rect 419172 22636 419224 22642
rect 419172 22578 419224 22584
rect 419184 17202 419212 22578
rect 419276 17542 419304 106286
rect 419264 17536 419316 17542
rect 419264 17478 419316 17484
rect 419736 17338 419764 107034
rect 419724 17332 419776 17338
rect 419724 17274 419776 17280
rect 419828 17270 419856 107102
rect 419920 106962 419948 456078
rect 419908 106956 419960 106962
rect 419908 106898 419960 106904
rect 419816 17264 419868 17270
rect 419816 17206 419868 17212
rect 419172 17196 419224 17202
rect 419172 17138 419224 17144
rect 419920 16454 419948 106898
rect 420012 106214 420040 479470
rect 436204 463146 436232 496975
rect 437492 496913 437520 497626
rect 438860 497616 438912 497622
rect 438860 497558 438912 497564
rect 438872 496913 438900 497558
rect 437478 496904 437534 496913
rect 437478 496839 437534 496848
rect 438858 496904 438914 496913
rect 438858 496839 438914 496848
rect 440238 496904 440294 496913
rect 440238 496839 440294 496848
rect 436192 463140 436244 463146
rect 436192 463082 436244 463088
rect 437492 456278 437520 496839
rect 437480 456272 437532 456278
rect 437480 456214 437532 456220
rect 438872 456210 438900 496839
rect 440252 465050 440280 496839
rect 441632 494057 441660 498063
rect 445312 497758 445340 498063
rect 445300 497752 445352 497758
rect 445300 497694 445352 497700
rect 444196 497684 444248 497690
rect 444196 497626 444248 497632
rect 444208 497457 444236 497626
rect 444194 497448 444250 497457
rect 444194 497383 444250 497392
rect 443644 497208 443696 497214
rect 443644 497150 443696 497156
rect 443656 496913 443684 497150
rect 443642 496904 443698 496913
rect 443642 496839 443698 496848
rect 441618 494048 441674 494057
rect 441618 493983 441674 493992
rect 443656 483886 443684 496839
rect 444208 494902 444236 497383
rect 444196 494896 444248 494902
rect 444196 494838 444248 494844
rect 445312 490686 445340 497694
rect 449176 497418 449204 498063
rect 451292 497554 451320 498063
rect 451280 497548 451332 497554
rect 451280 497490 451332 497496
rect 452396 497486 452424 498063
rect 452384 497480 452436 497486
rect 450542 497448 450598 497457
rect 449164 497412 449216 497418
rect 452384 497422 452436 497428
rect 450542 497383 450598 497392
rect 449164 497354 449216 497360
rect 447784 497276 447836 497282
rect 447784 497218 447836 497224
rect 446678 497176 446734 497185
rect 446678 497111 446734 497120
rect 446692 497078 446720 497111
rect 446680 497072 446732 497078
rect 447796 497049 447824 497218
rect 446680 497014 446732 497020
rect 447782 497040 447838 497049
rect 446692 496738 446720 497014
rect 447782 496975 447838 496984
rect 447138 496904 447194 496913
rect 447138 496839 447194 496848
rect 445760 496732 445812 496738
rect 445760 496674 445812 496680
rect 446680 496732 446732 496738
rect 446680 496674 446732 496680
rect 445300 490680 445352 490686
rect 445300 490622 445352 490628
rect 443644 483880 443696 483886
rect 443644 483822 443696 483828
rect 440240 465044 440292 465050
rect 440240 464986 440292 464992
rect 445772 463010 445800 496674
rect 447152 479670 447180 496839
rect 447140 479664 447192 479670
rect 447140 479606 447192 479612
rect 447796 469198 447824 496975
rect 449176 481642 449204 497354
rect 450556 497350 450584 497383
rect 450544 497344 450596 497350
rect 450544 497286 450596 497292
rect 449898 496904 449954 496913
rect 449898 496839 449954 496848
rect 449912 486674 449940 496839
rect 449900 486668 449952 486674
rect 449900 486610 449952 486616
rect 449164 481636 449216 481642
rect 449164 481578 449216 481584
rect 450556 470558 450584 497286
rect 453302 497040 453358 497049
rect 453302 496975 453358 496984
rect 453316 496942 453344 496975
rect 453304 496936 453356 496942
rect 452658 496904 452714 496913
rect 453304 496878 453356 496884
rect 452658 496839 452714 496848
rect 452672 489258 452700 496839
rect 452660 489252 452712 489258
rect 452660 489194 452712 489200
rect 453316 479534 453344 496878
rect 454604 489914 454632 498063
rect 454604 489886 454724 489914
rect 453304 479528 453356 479534
rect 453304 479470 453356 479476
rect 450544 470552 450596 470558
rect 450544 470494 450596 470500
rect 447784 469192 447836 469198
rect 447784 469134 447836 469140
rect 445760 463004 445812 463010
rect 445760 462946 445812 462952
rect 438860 456204 438912 456210
rect 438860 456146 438912 456152
rect 454696 456142 454724 489886
rect 455524 488034 455552 498063
rect 463698 497992 463754 498001
rect 463698 497927 463754 497936
rect 467838 497992 467894 498001
rect 467838 497927 467894 497936
rect 460570 497856 460626 497865
rect 460570 497791 460626 497800
rect 462318 497856 462374 497865
rect 462318 497791 462374 497800
rect 457442 497448 457498 497457
rect 457442 497383 457498 497392
rect 456064 497140 456116 497146
rect 456064 497082 456116 497088
rect 456076 496913 456104 497082
rect 456062 496904 456118 496913
rect 456062 496839 456118 496848
rect 456890 496904 456946 496913
rect 456890 496839 456946 496848
rect 456076 488510 456104 496839
rect 456904 492658 456932 496839
rect 456892 492652 456944 492658
rect 456892 492594 456944 492600
rect 456064 488504 456116 488510
rect 456064 488446 456116 488452
rect 455512 488028 455564 488034
rect 455512 487970 455564 487976
rect 457456 471986 457484 497383
rect 460584 497010 460612 497791
rect 462332 497690 462360 497791
rect 463712 497758 463740 497927
rect 463700 497752 463752 497758
rect 463700 497694 463752 497700
rect 462320 497684 462372 497690
rect 462320 497626 462372 497632
rect 462504 497684 462556 497690
rect 462504 497626 462556 497632
rect 462044 497616 462096 497622
rect 462044 497558 462096 497564
rect 461122 497312 461178 497321
rect 461122 497247 461178 497256
rect 461136 497214 461164 497247
rect 461124 497208 461176 497214
rect 461124 497150 461176 497156
rect 462056 497049 462084 497558
rect 462516 497457 462544 497626
rect 462502 497448 462558 497457
rect 462502 497383 462558 497392
rect 466458 497448 466514 497457
rect 466458 497383 466460 497392
rect 466512 497383 466514 497392
rect 466460 497354 466512 497360
rect 467852 497350 467880 497927
rect 469232 497554 469260 498063
rect 470874 497720 470930 497729
rect 470874 497655 470930 497664
rect 469220 497548 469272 497554
rect 469220 497490 469272 497496
rect 470888 497486 470916 497655
rect 470876 497480 470928 497486
rect 470876 497422 470928 497428
rect 467840 497344 467892 497350
rect 465078 497312 465134 497321
rect 467840 497286 467892 497292
rect 465078 497247 465080 497256
rect 465132 497247 465134 497256
rect 465080 497218 465132 497224
rect 465078 497176 465134 497185
rect 465078 497111 465134 497120
rect 473358 497176 473414 497185
rect 473358 497111 473360 497120
rect 465092 497078 465120 497111
rect 473412 497111 473414 497120
rect 473360 497082 473412 497088
rect 465080 497072 465132 497078
rect 462042 497040 462098 497049
rect 459560 497004 459612 497010
rect 459560 496946 459612 496952
rect 460572 497004 460624 497010
rect 465080 497014 465132 497020
rect 471978 497040 472034 497049
rect 462042 496975 462098 496984
rect 471978 496975 472034 496984
rect 460572 496946 460624 496952
rect 458178 496904 458234 496913
rect 459466 496904 459522 496913
rect 458178 496839 458234 496848
rect 458824 496868 458876 496874
rect 458192 483818 458220 496839
rect 459466 496839 459468 496848
rect 458824 496810 458876 496816
rect 459520 496839 459522 496848
rect 459468 496810 459520 496816
rect 458180 483812 458232 483818
rect 458180 483754 458232 483760
rect 457444 471980 457496 471986
rect 457444 471922 457496 471928
rect 458836 466410 458864 496810
rect 459572 496806 459600 496946
rect 471992 496942 472020 496975
rect 471980 496936 472032 496942
rect 460938 496904 460994 496913
rect 460938 496839 460994 496848
rect 462410 496904 462466 496913
rect 462410 496839 462466 496848
rect 465170 496904 465226 496913
rect 465170 496839 465226 496848
rect 467930 496904 467986 496913
rect 467930 496839 467986 496848
rect 470782 496904 470838 496913
rect 471980 496878 472032 496884
rect 470782 496839 470838 496848
rect 459560 496800 459612 496806
rect 459560 496742 459612 496748
rect 460952 490754 460980 496839
rect 460940 490748 460992 490754
rect 460940 490690 460992 490696
rect 462424 482526 462452 496839
rect 462412 482520 462464 482526
rect 462412 482462 462464 482468
rect 465184 481098 465212 496839
rect 465172 481092 465224 481098
rect 465172 481034 465224 481040
rect 467944 471306 467972 496839
rect 470796 496126 470824 496839
rect 470784 496120 470836 496126
rect 470784 496062 470836 496068
rect 473556 494834 473584 498063
rect 474738 497720 474794 497729
rect 474738 497655 474794 497664
rect 476118 497720 476174 497729
rect 476118 497655 476120 497664
rect 474752 497622 474780 497655
rect 476172 497655 476174 497664
rect 476120 497626 476172 497632
rect 474740 497616 474792 497622
rect 474740 497558 474792 497564
rect 478878 497312 478934 497321
rect 478878 497247 478934 497256
rect 477590 497040 477646 497049
rect 478892 497010 478920 497247
rect 477590 496975 477646 496984
rect 478880 497004 478932 497010
rect 476118 496904 476174 496913
rect 476118 496839 476174 496848
rect 477498 496904 477554 496913
rect 477498 496839 477500 496848
rect 473544 494828 473596 494834
rect 473544 494770 473596 494776
rect 476132 476814 476160 496839
rect 477552 496839 477554 496848
rect 477500 496810 477552 496816
rect 477604 493474 477632 496975
rect 478880 496946 478932 496952
rect 477592 493468 477644 493474
rect 477592 493410 477644 493416
rect 480548 492046 480576 498063
rect 483018 496904 483074 496913
rect 483018 496839 483074 496848
rect 485778 496904 485834 496913
rect 485778 496839 485834 496848
rect 487158 496904 487214 496913
rect 487158 496839 487214 496848
rect 490470 496904 490526 496913
rect 490470 496839 490526 496848
rect 492678 496904 492734 496913
rect 492678 496839 492734 496848
rect 480536 492040 480588 492046
rect 480536 491982 480588 491988
rect 483032 478242 483060 496839
rect 485792 480962 485820 496839
rect 487172 482390 487200 496839
rect 490484 490618 490512 496839
rect 490472 490612 490524 490618
rect 490472 490554 490524 490560
rect 492692 483750 492720 496839
rect 492680 483744 492732 483750
rect 492680 483686 492732 483692
rect 487160 482384 487212 482390
rect 487160 482326 487212 482332
rect 485780 480956 485832 480962
rect 485780 480898 485832 480904
rect 483020 478236 483072 478242
rect 483020 478178 483072 478184
rect 476120 476808 476172 476814
rect 476120 476750 476172 476756
rect 467932 471300 467984 471306
rect 467932 471242 467984 471248
rect 458824 466404 458876 466410
rect 458824 466346 458876 466352
rect 494716 461650 494744 498063
rect 497462 496904 497518 496913
rect 497462 496839 497518 496848
rect 500958 496904 501014 496913
rect 500958 496839 501014 496848
rect 502338 496904 502394 496913
rect 502338 496839 502394 496848
rect 497476 487830 497504 496839
rect 500972 489190 501000 496839
rect 500960 489184 501012 489190
rect 500960 489126 501012 489132
rect 497464 487824 497516 487830
rect 497464 487766 497516 487772
rect 502352 475386 502380 496839
rect 502340 475380 502392 475386
rect 502340 475322 502392 475328
rect 504376 472666 504404 498063
rect 507858 496904 507914 496913
rect 507858 496839 507914 496848
rect 510618 496904 510674 496913
rect 510618 496839 510674 496848
rect 504364 472660 504416 472666
rect 504364 472602 504416 472608
rect 507872 468518 507900 496839
rect 507860 468512 507912 468518
rect 507860 468454 507912 468460
rect 510632 465798 510660 496839
rect 512656 467158 512684 498063
rect 514758 496904 514814 496913
rect 514758 496839 514814 496848
rect 517518 496904 517574 496913
rect 517518 496839 517574 496848
rect 514772 469878 514800 496839
rect 514760 469872 514812 469878
rect 514760 469814 514812 469820
rect 512644 467152 512696 467158
rect 512644 467094 512696 467100
rect 510620 465792 510672 465798
rect 510620 465734 510672 465740
rect 517532 464438 517560 496839
rect 517520 464432 517572 464438
rect 517520 464374 517572 464380
rect 519556 463078 519584 498063
rect 523038 496904 523094 496913
rect 523038 496839 523094 496848
rect 525798 496904 525854 496913
rect 525798 496839 525854 496848
rect 523052 474094 523080 496839
rect 523040 474088 523092 474094
rect 523040 474030 523092 474036
rect 519544 463072 519596 463078
rect 519544 463014 519596 463020
rect 494704 461644 494756 461650
rect 494704 461586 494756 461592
rect 454684 456136 454736 456142
rect 454684 456078 454736 456084
rect 525812 454714 525840 496839
rect 558288 474026 558316 510614
rect 558276 474020 558328 474026
rect 558276 473962 558328 473968
rect 525800 454708 525852 454714
rect 525800 454650 525852 454656
rect 558182 454200 558238 454209
rect 558182 454135 558238 454144
rect 551006 196072 551062 196081
rect 551006 196007 551008 196016
rect 551060 196007 551062 196016
rect 557540 196036 557592 196042
rect 551008 195978 551060 195984
rect 557540 195978 557592 195984
rect 451278 109848 451334 109857
rect 451278 109783 451334 109792
rect 480902 109848 480958 109857
rect 480902 109783 480958 109792
rect 483478 109848 483534 109857
rect 483478 109783 483534 109792
rect 485962 109848 486018 109857
rect 485962 109783 486018 109792
rect 488262 109848 488318 109857
rect 488262 109783 488318 109792
rect 491022 109848 491078 109857
rect 491022 109783 491078 109792
rect 451292 109750 451320 109783
rect 451280 109744 451332 109750
rect 451280 109686 451332 109692
rect 452476 109744 452528 109750
rect 452476 109686 452528 109692
rect 476118 109712 476174 109721
rect 450636 107636 450688 107642
rect 450636 107578 450688 107584
rect 450648 107545 450676 107578
rect 436098 107536 436154 107545
rect 436098 107471 436154 107480
rect 437018 107536 437074 107545
rect 437018 107471 437074 107480
rect 438122 107536 438178 107545
rect 438122 107471 438178 107480
rect 439594 107536 439650 107545
rect 439594 107471 439650 107480
rect 440514 107536 440570 107545
rect 440514 107471 440570 107480
rect 441618 107536 441674 107545
rect 441618 107471 441674 107480
rect 443090 107536 443146 107545
rect 443090 107471 443146 107480
rect 444194 107536 444250 107545
rect 444194 107471 444250 107480
rect 445666 107536 445722 107545
rect 445666 107471 445722 107480
rect 446402 107536 446458 107545
rect 446402 107471 446458 107480
rect 447138 107536 447194 107545
rect 447138 107471 447194 107480
rect 448518 107536 448574 107545
rect 448518 107471 448574 107480
rect 449898 107536 449954 107545
rect 449898 107471 449954 107480
rect 450634 107536 450690 107545
rect 450634 107471 450690 107480
rect 436112 107234 436140 107471
rect 436100 107228 436152 107234
rect 436100 107170 436152 107176
rect 437032 106894 437060 107471
rect 438136 107166 438164 107471
rect 438124 107160 438176 107166
rect 438124 107102 438176 107108
rect 439608 107098 439636 107471
rect 439596 107092 439648 107098
rect 439596 107034 439648 107040
rect 437020 106888 437072 106894
rect 437020 106830 437072 106836
rect 440528 106486 440556 107471
rect 440516 106480 440568 106486
rect 440516 106422 440568 106428
rect 441632 106418 441660 107471
rect 441620 106412 441672 106418
rect 441620 106354 441672 106360
rect 443104 106350 443132 107471
rect 444208 107098 444236 107471
rect 444288 107160 444340 107166
rect 444288 107102 444340 107108
rect 444196 107092 444248 107098
rect 444196 107034 444248 107040
rect 444300 106350 444328 107102
rect 445680 106486 445708 107471
rect 445668 106480 445720 106486
rect 445668 106422 445720 106428
rect 443092 106344 443144 106350
rect 443092 106286 443144 106292
rect 444288 106344 444340 106350
rect 444288 106286 444340 106292
rect 420000 106208 420052 106214
rect 420000 106150 420052 106156
rect 419908 16448 419960 16454
rect 419908 16390 419960 16396
rect 420012 16318 420040 106150
rect 445680 106010 445708 106422
rect 446416 106418 446444 107471
rect 447152 106622 447180 107471
rect 448532 106690 448560 107471
rect 448520 106684 448572 106690
rect 448520 106626 448572 106632
rect 447140 106616 447192 106622
rect 447140 106558 447192 106564
rect 446404 106412 446456 106418
rect 446404 106354 446456 106360
rect 446416 106078 446444 106354
rect 447152 106146 447180 106558
rect 447140 106140 447192 106146
rect 447140 106082 447192 106088
rect 446404 106072 446456 106078
rect 446404 106014 446456 106020
rect 445668 106004 445720 106010
rect 445668 105946 445720 105952
rect 448532 105602 448560 106626
rect 449912 106554 449940 107471
rect 452488 107302 452516 109686
rect 480916 109682 480944 109783
rect 476118 109647 476174 109656
rect 480904 109676 480956 109682
rect 456982 109576 457038 109585
rect 456982 109511 457038 109520
rect 452568 107976 452620 107982
rect 452568 107918 452620 107924
rect 452580 107545 452608 107918
rect 456996 107914 457024 109511
rect 476132 109138 476160 109647
rect 480904 109618 480956 109624
rect 483492 109614 483520 109783
rect 483480 109608 483532 109614
rect 483480 109550 483532 109556
rect 485976 109546 486004 109783
rect 485964 109540 486016 109546
rect 485964 109482 486016 109488
rect 488276 109478 488304 109783
rect 488264 109472 488316 109478
rect 488264 109414 488316 109420
rect 491036 109410 491064 109783
rect 493414 109712 493470 109721
rect 493414 109647 493470 109656
rect 495898 109712 495954 109721
rect 495898 109647 495954 109656
rect 498474 109712 498530 109721
rect 498474 109647 498530 109656
rect 491024 109404 491076 109410
rect 491024 109346 491076 109352
rect 493428 109342 493456 109647
rect 493416 109336 493468 109342
rect 493416 109278 493468 109284
rect 495912 109274 495940 109647
rect 495900 109268 495952 109274
rect 495900 109210 495952 109216
rect 498488 109206 498516 109647
rect 505926 109576 505982 109585
rect 505926 109511 505982 109520
rect 508502 109576 508558 109585
rect 508502 109511 508558 109520
rect 515862 109576 515918 109585
rect 515862 109511 515918 109520
rect 518438 109576 518494 109585
rect 518438 109511 518494 109520
rect 498476 109200 498528 109206
rect 498476 109142 498528 109148
rect 476120 109132 476172 109138
rect 476120 109074 476172 109080
rect 500958 109032 501014 109041
rect 500958 108967 501014 108976
rect 503442 109032 503498 109041
rect 503442 108967 503498 108976
rect 500972 108866 501000 108967
rect 500960 108860 501012 108866
rect 500960 108802 501012 108808
rect 503456 108798 503484 108967
rect 503444 108792 503496 108798
rect 503444 108734 503496 108740
rect 505940 108730 505968 109511
rect 508516 109070 508544 109511
rect 508504 109064 508556 109070
rect 508504 109006 508556 109012
rect 513378 109032 513434 109041
rect 513378 108967 513434 108976
rect 505928 108724 505980 108730
rect 505928 108666 505980 108672
rect 513392 108594 513420 108967
rect 513380 108588 513432 108594
rect 513380 108530 513432 108536
rect 515876 108526 515904 109511
rect 515864 108520 515916 108526
rect 457994 108488 458050 108497
rect 515864 108462 515916 108468
rect 518452 108458 518480 109511
rect 520922 109032 520978 109041
rect 520922 108967 520978 108976
rect 523314 109032 523370 109041
rect 523314 108967 523370 108976
rect 525890 109032 525946 109041
rect 525890 108967 525946 108976
rect 520936 108662 520964 108967
rect 520924 108656 520976 108662
rect 520924 108598 520976 108604
rect 457994 108423 458050 108432
rect 518440 108452 518492 108458
rect 458008 108050 458036 108423
rect 518440 108394 518492 108400
rect 523328 108322 523356 108967
rect 525904 108390 525932 108967
rect 525892 108384 525944 108390
rect 525892 108326 525944 108332
rect 523316 108316 523368 108322
rect 523316 108258 523368 108264
rect 457996 108044 458048 108050
rect 457996 107986 458048 107992
rect 456984 107908 457036 107914
rect 456984 107850 457036 107856
rect 455788 107840 455840 107846
rect 455788 107782 455840 107788
rect 455800 107545 455828 107782
rect 456996 107710 457024 107850
rect 456984 107704 457036 107710
rect 456984 107646 457036 107652
rect 452566 107536 452622 107545
rect 452566 107471 452622 107480
rect 453578 107536 453634 107545
rect 453578 107471 453634 107480
rect 454590 107536 454646 107545
rect 454590 107471 454646 107480
rect 455786 107536 455842 107545
rect 455786 107471 455842 107480
rect 455970 107536 456026 107545
rect 455970 107471 455972 107480
rect 452580 107370 452608 107471
rect 452568 107364 452620 107370
rect 452568 107306 452620 107312
rect 452476 107296 452528 107302
rect 452476 107238 452528 107244
rect 453592 106826 453620 107471
rect 453946 107128 454002 107137
rect 453946 107063 454002 107072
rect 453580 106820 453632 106826
rect 453580 106762 453632 106768
rect 449900 106548 449952 106554
rect 449900 106490 449952 106496
rect 449912 105670 449940 106490
rect 453960 106350 453988 107063
rect 454604 107030 454632 107471
rect 455800 107438 455828 107471
rect 456024 107471 456026 107480
rect 455972 107442 456024 107448
rect 455788 107432 455840 107438
rect 455788 107374 455840 107380
rect 458008 107137 458036 107986
rect 458180 107772 458232 107778
rect 458180 107714 458232 107720
rect 458192 107642 458220 107714
rect 458180 107636 458232 107642
rect 458180 107578 458232 107584
rect 459468 107636 459520 107642
rect 459468 107578 459520 107584
rect 475660 107636 475712 107642
rect 475660 107578 475712 107584
rect 458364 107568 458416 107574
rect 458362 107536 458364 107545
rect 459480 107545 459508 107578
rect 475672 107545 475700 107578
rect 478052 107568 478104 107574
rect 458416 107536 458418 107545
rect 458362 107471 458418 107480
rect 459466 107536 459522 107545
rect 459466 107471 459522 107480
rect 460662 107536 460718 107545
rect 460662 107471 460718 107480
rect 461674 107536 461730 107545
rect 461674 107471 461730 107480
rect 462778 107536 462834 107545
rect 462778 107471 462834 107480
rect 463882 107536 463938 107545
rect 463882 107471 463938 107480
rect 465170 107536 465226 107545
rect 465170 107471 465226 107480
rect 465722 107536 465778 107545
rect 465722 107471 465778 107480
rect 467010 107536 467066 107545
rect 467010 107471 467066 107480
rect 468666 107536 468722 107545
rect 468666 107471 468722 107480
rect 469770 107536 469826 107545
rect 469770 107471 469826 107480
rect 471150 107536 471206 107545
rect 471150 107471 471206 107480
rect 472070 107536 472126 107545
rect 472070 107471 472126 107480
rect 473358 107536 473414 107545
rect 473358 107471 473414 107480
rect 474370 107536 474426 107545
rect 474370 107471 474372 107480
rect 459560 107228 459612 107234
rect 459560 107170 459612 107176
rect 457994 107128 458050 107137
rect 457994 107063 458050 107072
rect 454592 107024 454644 107030
rect 454592 106966 454644 106972
rect 459572 106962 459600 107170
rect 460676 106962 460704 107471
rect 461688 107166 461716 107471
rect 461676 107160 461728 107166
rect 461676 107102 461728 107108
rect 462792 107098 462820 107471
rect 462780 107092 462832 107098
rect 462780 107034 462832 107040
rect 459560 106956 459612 106962
rect 459560 106898 459612 106904
rect 460664 106956 460716 106962
rect 460664 106898 460716 106904
rect 463896 106486 463924 107471
rect 463884 106480 463936 106486
rect 463884 106422 463936 106428
rect 465184 106418 465212 107471
rect 465736 106622 465764 107471
rect 467024 106690 467052 107471
rect 467012 106684 467064 106690
rect 467012 106626 467064 106632
rect 465724 106616 465776 106622
rect 465724 106558 465776 106564
rect 468680 106554 468708 107471
rect 469784 107302 469812 107471
rect 471164 107438 471192 107471
rect 471152 107432 471204 107438
rect 471152 107374 471204 107380
rect 469772 107296 469824 107302
rect 469772 107238 469824 107244
rect 468668 106548 468720 106554
rect 468668 106490 468720 106496
rect 465172 106412 465224 106418
rect 465172 106354 465224 106360
rect 472084 106350 472112 107471
rect 473372 107030 473400 107471
rect 474424 107471 474426 107480
rect 475658 107536 475714 107545
rect 475658 107471 475714 107480
rect 478050 107536 478052 107545
rect 478104 107536 478106 107545
rect 478050 107471 478106 107480
rect 479154 107536 479210 107545
rect 479154 107471 479210 107480
rect 474372 107442 474424 107448
rect 473360 107024 473412 107030
rect 473360 106966 473412 106972
rect 479168 106962 479196 107471
rect 479156 106956 479208 106962
rect 479156 106898 479208 106904
rect 453948 106344 454000 106350
rect 453948 106286 454000 106292
rect 472072 106344 472124 106350
rect 472072 106286 472124 106292
rect 453960 106214 453988 106286
rect 557552 106282 557580 195978
rect 550732 106276 550784 106282
rect 550732 106218 550784 106224
rect 557540 106276 557592 106282
rect 557540 106218 557592 106224
rect 453948 106208 454000 106214
rect 453948 106150 454000 106156
rect 449900 105664 449952 105670
rect 449900 105606 449952 105612
rect 448520 105596 448572 105602
rect 448520 105538 448572 105544
rect 550744 105369 550772 106218
rect 550730 105360 550786 105369
rect 550730 105295 550786 105304
rect 558196 46918 558224 454135
rect 558932 247790 558960 579119
rect 562324 563100 562376 563106
rect 562324 563042 562376 563048
rect 562336 478174 562364 563042
rect 562324 478168 562376 478174
rect 562324 478110 562376 478116
rect 563716 457502 563744 616830
rect 565096 457570 565124 670686
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 569224 643136 569276 643142
rect 569224 643078 569276 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 566464 536852 566516 536858
rect 566464 536794 566516 536800
rect 566476 482322 566504 536794
rect 569236 493338 569264 643078
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 573364 630692 573416 630698
rect 573364 630634 573416 630640
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 571984 576904 572036 576910
rect 571984 576846 572036 576852
rect 570604 524476 570656 524482
rect 570604 524418 570656 524424
rect 569224 493332 569276 493338
rect 569224 493274 569276 493280
rect 570616 483682 570644 524418
rect 571996 494766 572024 576846
rect 571984 494760 572036 494766
rect 571984 494702 572036 494708
rect 573376 486470 573404 630634
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 573364 486464 573416 486470
rect 573364 486406 573416 486412
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 570604 483676 570656 483682
rect 570604 483618 570656 483624
rect 566464 482316 566516 482322
rect 566464 482258 566516 482264
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580632 460964 580684 460970
rect 580632 460906 580684 460912
rect 580538 458416 580594 458425
rect 580538 458351 580594 458360
rect 580448 458312 580500 458318
rect 580354 458280 580410 458289
rect 580448 458254 580500 458260
rect 580354 458215 580410 458224
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 565084 457564 565136 457570
rect 565084 457506 565136 457512
rect 563704 457496 563756 457502
rect 563704 457438 563756 457444
rect 580184 456074 580212 458079
rect 580172 456068 580224 456074
rect 580172 456010 580224 456016
rect 573362 455696 573418 455705
rect 573362 455631 573418 455640
rect 571982 455560 572038 455569
rect 571982 455495 572038 455504
rect 562324 455456 562376 455462
rect 562324 455398 562376 455404
rect 558920 247784 558972 247790
rect 558920 247726 558972 247732
rect 558932 189145 558960 247726
rect 562336 193186 562364 455398
rect 570604 454096 570656 454102
rect 566462 454064 566518 454073
rect 570604 454038 570656 454044
rect 566462 453999 566518 454008
rect 565820 243568 565872 243574
rect 565820 243510 565872 243516
rect 565084 242208 565136 242214
rect 565084 242150 565136 242156
rect 562416 199436 562468 199442
rect 562416 199378 562468 199384
rect 562324 193180 562376 193186
rect 562324 193122 562376 193128
rect 558918 189136 558974 189145
rect 558918 189071 558974 189080
rect 558932 99385 558960 189071
rect 558918 99376 558974 99385
rect 558918 99311 558974 99320
rect 558184 46912 558236 46918
rect 558184 46854 558236 46860
rect 460662 19816 460718 19825
rect 460662 19751 460664 19760
rect 460716 19751 460718 19760
rect 488262 19816 488318 19825
rect 488262 19751 488318 19760
rect 460664 19722 460716 19728
rect 447598 19680 447654 19689
rect 447598 19615 447654 19624
rect 448702 19680 448758 19689
rect 448702 19615 448758 19624
rect 450082 19680 450138 19689
rect 450082 19615 450138 19624
rect 455970 19680 456026 19689
rect 455970 19615 456026 19624
rect 447612 19310 447640 19615
rect 447600 19304 447652 19310
rect 447600 19246 447652 19252
rect 445668 18488 445720 18494
rect 445668 18430 445720 18436
rect 444288 18420 444340 18426
rect 444288 18362 444340 18368
rect 444300 17921 444328 18362
rect 445680 17921 445708 18430
rect 436098 17912 436154 17921
rect 436098 17847 436154 17856
rect 436282 17912 436338 17921
rect 436282 17847 436338 17856
rect 437478 17912 437534 17921
rect 437478 17847 437534 17856
rect 438858 17912 438914 17921
rect 438858 17847 438914 17856
rect 440238 17912 440294 17921
rect 440238 17847 440294 17856
rect 441710 17912 441766 17921
rect 441710 17847 441766 17856
rect 443090 17912 443146 17921
rect 443090 17847 443146 17856
rect 444286 17912 444342 17921
rect 444286 17847 444288 17856
rect 436112 17202 436140 17847
rect 436100 17196 436152 17202
rect 436100 17138 436152 17144
rect 436296 17134 436324 17847
rect 437492 17270 437520 17847
rect 438872 17338 438900 17847
rect 440252 17406 440280 17847
rect 441724 17474 441752 17847
rect 443104 17542 443132 17847
rect 444340 17847 444342 17856
rect 445666 17912 445722 17921
rect 445666 17847 445722 17856
rect 446494 17912 446550 17921
rect 446494 17847 446550 17856
rect 447138 17912 447194 17921
rect 447138 17847 447194 17856
rect 444288 17818 444340 17824
rect 444300 17787 444328 17818
rect 445680 17678 445708 17847
rect 445668 17672 445720 17678
rect 445668 17614 445720 17620
rect 443092 17536 443144 17542
rect 443092 17478 443144 17484
rect 441712 17468 441764 17474
rect 441712 17410 441764 17416
rect 440240 17400 440292 17406
rect 440240 17342 440292 17348
rect 438860 17332 438912 17338
rect 438860 17274 438912 17280
rect 437480 17264 437532 17270
rect 437480 17206 437532 17212
rect 436284 17128 436336 17134
rect 436284 17070 436336 17076
rect 446508 16998 446536 17847
rect 447152 17066 447180 17847
rect 447612 17474 447640 19246
rect 448716 19242 448744 19615
rect 448704 19236 448756 19242
rect 448704 19178 448756 19184
rect 448716 17610 448744 19178
rect 450096 18562 450124 19615
rect 455984 19174 456012 19615
rect 455972 19168 456024 19174
rect 455972 19110 456024 19116
rect 450084 18556 450136 18562
rect 450084 18498 450136 18504
rect 449898 17912 449954 17921
rect 449898 17847 449954 17856
rect 448704 17604 448756 17610
rect 448704 17546 448756 17552
rect 447600 17468 447652 17474
rect 447600 17410 447652 17416
rect 447140 17060 447192 17066
rect 447140 17002 447192 17008
rect 446496 16992 446548 16998
rect 446496 16934 446548 16940
rect 449912 16930 449940 17847
rect 450096 17542 450124 18498
rect 451278 17912 451334 17921
rect 451278 17847 451334 17856
rect 452290 17912 452346 17921
rect 452290 17847 452346 17856
rect 453486 17912 453542 17921
rect 453486 17847 453542 17856
rect 454038 17912 454094 17921
rect 454038 17847 454094 17856
rect 455418 17912 455474 17921
rect 455418 17847 455474 17856
rect 450084 17536 450136 17542
rect 450084 17478 450136 17484
rect 451292 16930 451320 17847
rect 449900 16924 449952 16930
rect 449900 16866 449952 16872
rect 451280 16924 451332 16930
rect 451280 16866 451332 16872
rect 451292 16386 451320 16866
rect 452304 16794 452332 17847
rect 451372 16788 451424 16794
rect 451372 16730 451424 16736
rect 452292 16788 452344 16794
rect 452292 16730 452344 16736
rect 451280 16380 451332 16386
rect 451280 16322 451332 16328
rect 420000 16312 420052 16318
rect 420000 16254 420052 16260
rect 451384 16250 451412 16730
rect 453500 16726 453528 17847
rect 452660 16720 452712 16726
rect 452660 16662 452712 16668
rect 453488 16720 453540 16726
rect 453488 16662 453540 16668
rect 452672 16318 452700 16662
rect 454052 16454 454080 17847
rect 455432 17814 455460 17847
rect 455984 17814 456012 19110
rect 458362 18048 458418 18057
rect 458362 17983 458418 17992
rect 458376 17950 458404 17983
rect 460676 17950 460704 19722
rect 488276 19718 488304 19751
rect 488264 19712 488316 19718
rect 473358 19680 473414 19689
rect 473414 19638 473492 19666
rect 488264 19654 488316 19660
rect 491022 19680 491078 19689
rect 473358 19615 473414 19624
rect 468298 19544 468354 19553
rect 468298 19479 468354 19488
rect 468312 19106 468340 19479
rect 468300 19100 468352 19106
rect 468300 19042 468352 19048
rect 470876 19032 470928 19038
rect 470876 18974 470928 18980
rect 470888 18873 470916 18974
rect 470874 18864 470930 18873
rect 470874 18799 470930 18808
rect 458364 17944 458416 17950
rect 457350 17912 457406 17921
rect 457350 17847 457406 17856
rect 458086 17912 458142 17921
rect 458086 17847 458142 17856
rect 458270 17912 458326 17921
rect 460664 17944 460716 17950
rect 458364 17886 458416 17892
rect 459466 17912 459522 17921
rect 458270 17847 458326 17856
rect 460664 17886 460716 17892
rect 462318 17912 462374 17921
rect 459466 17847 459522 17856
rect 462318 17847 462320 17856
rect 455420 17808 455472 17814
rect 455420 17750 455472 17756
rect 455972 17808 456024 17814
rect 455972 17750 456024 17756
rect 456800 17740 456852 17746
rect 456800 17682 456852 17688
rect 456812 17338 456840 17682
rect 456800 17332 456852 17338
rect 456800 17274 456852 17280
rect 457364 16862 457392 17847
rect 458100 17338 458128 17847
rect 458088 17332 458140 17338
rect 458088 17274 458140 17280
rect 457352 16856 457404 16862
rect 457352 16798 457404 16804
rect 457364 16522 457392 16798
rect 458284 16590 458312 17847
rect 459480 17406 459508 17847
rect 462372 17847 462374 17856
rect 463698 17912 463754 17921
rect 463698 17847 463754 17856
rect 465078 17912 465134 17921
rect 465078 17847 465134 17856
rect 466458 17912 466514 17921
rect 466458 17847 466514 17856
rect 467838 17912 467894 17921
rect 467838 17847 467894 17856
rect 473358 17912 473414 17921
rect 473358 17847 473414 17856
rect 462320 17818 462372 17824
rect 463712 17678 463740 17847
rect 463700 17672 463752 17678
rect 463700 17614 463752 17620
rect 465092 17474 465120 17847
rect 466472 17610 466500 17847
rect 466460 17604 466512 17610
rect 466460 17546 466512 17552
rect 467852 17542 467880 17847
rect 473372 17814 473400 17847
rect 473360 17808 473412 17814
rect 473360 17750 473412 17756
rect 467840 17536 467892 17542
rect 467840 17478 467892 17484
rect 465080 17468 465132 17474
rect 465080 17410 465132 17416
rect 459468 17400 459520 17406
rect 459468 17342 459520 17348
rect 471702 17368 471758 17377
rect 471702 17303 471758 17312
rect 465080 17264 465132 17270
rect 465080 17206 465132 17212
rect 465092 17105 465120 17206
rect 471716 17105 471744 17303
rect 471978 17232 472034 17241
rect 471978 17167 472034 17176
rect 465078 17096 465134 17105
rect 465078 17031 465134 17040
rect 469310 17096 469366 17105
rect 469310 17031 469366 17040
rect 471702 17096 471758 17105
rect 471702 17031 471758 17040
rect 469324 16998 469352 17031
rect 469312 16992 469364 16998
rect 469312 16934 469364 16940
rect 469220 16924 469272 16930
rect 469220 16866 469272 16872
rect 458272 16584 458324 16590
rect 458272 16526 458324 16532
rect 457352 16516 457404 16522
rect 457352 16458 457404 16464
rect 469232 16454 469260 16866
rect 470874 16824 470930 16833
rect 470874 16759 470876 16768
rect 470928 16759 470930 16768
rect 470876 16730 470928 16736
rect 471992 16726 472020 17167
rect 473464 16930 473492 19638
rect 491022 19615 491024 19624
rect 491076 19615 491078 19624
rect 493414 19680 493470 19689
rect 493414 19615 493470 19624
rect 491024 19586 491076 19592
rect 493428 19582 493456 19615
rect 493416 19576 493468 19582
rect 493416 19518 493468 19524
rect 495898 19544 495954 19553
rect 495898 19479 495900 19488
rect 495952 19479 495954 19488
rect 500958 19544 501014 19553
rect 500958 19479 501014 19488
rect 503534 19544 503590 19553
rect 503534 19479 503590 19488
rect 495900 19450 495952 19456
rect 500972 19446 501000 19479
rect 500960 19440 501012 19446
rect 500960 19382 501012 19388
rect 503548 19378 503576 19479
rect 503536 19372 503588 19378
rect 503536 19314 503588 19320
rect 485042 19272 485098 19281
rect 485042 19207 485098 19216
rect 498474 19272 498530 19281
rect 498474 19207 498530 19216
rect 501050 19272 501106 19281
rect 501050 19207 501106 19216
rect 485056 18873 485084 19207
rect 485042 18864 485098 18873
rect 485042 18799 485098 18808
rect 498488 18766 498516 19207
rect 501064 18873 501092 19207
rect 515770 19000 515826 19009
rect 515770 18935 515772 18944
rect 515824 18935 515826 18944
rect 515772 18906 515824 18912
rect 505836 18896 505888 18902
rect 501050 18864 501106 18873
rect 501050 18799 501106 18808
rect 505834 18864 505836 18873
rect 505888 18864 505890 18873
rect 505834 18799 505890 18808
rect 508410 18864 508466 18873
rect 508410 18799 508412 18808
rect 508464 18799 508466 18808
rect 508412 18770 508464 18776
rect 498476 18760 498528 18766
rect 498476 18702 498528 18708
rect 523314 18728 523370 18737
rect 523314 18663 523316 18672
rect 523368 18663 523370 18672
rect 525890 18728 525946 18737
rect 525890 18663 525946 18672
rect 523316 18634 523368 18640
rect 525904 18630 525932 18663
rect 525892 18624 525944 18630
rect 525892 18566 525944 18572
rect 478880 17944 478932 17950
rect 476118 17912 476174 17921
rect 476118 17847 476174 17856
rect 478878 17912 478880 17921
rect 478932 17912 478934 17921
rect 478878 17847 478934 17856
rect 475382 17776 475438 17785
rect 475382 17711 475438 17720
rect 475396 17513 475424 17711
rect 475382 17504 475438 17513
rect 475382 17439 475438 17448
rect 476132 17338 476160 17847
rect 476120 17332 476172 17338
rect 476120 17274 476172 17280
rect 474738 17232 474794 17241
rect 474738 17167 474794 17176
rect 473452 16924 473504 16930
rect 473452 16866 473504 16872
rect 474752 16862 474780 17167
rect 477498 16960 477554 16969
rect 477498 16895 477554 16904
rect 474740 16856 474792 16862
rect 474740 16798 474792 16804
rect 471980 16720 472032 16726
rect 471980 16662 472032 16668
rect 477512 16658 477540 16895
rect 477500 16652 477552 16658
rect 477500 16594 477552 16600
rect 454040 16448 454092 16454
rect 454040 16390 454092 16396
rect 469220 16448 469272 16454
rect 469220 16390 469272 16396
rect 452660 16312 452712 16318
rect 452660 16254 452712 16260
rect 451372 16244 451424 16250
rect 451372 16186 451424 16192
rect 420920 15972 420972 15978
rect 420920 15914 420972 15920
rect 419080 3324 419132 3330
rect 419080 3266 419132 3272
rect 418528 3256 418580 3262
rect 418528 3198 418580 3204
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 15914
rect 432052 15904 432104 15910
rect 432052 15846 432104 15852
rect 423680 14544 423732 14550
rect 423680 14486 423732 14492
rect 423692 3194 423720 14486
rect 428464 11824 428516 11830
rect 428464 11766 428516 11772
rect 423680 3188 423732 3194
rect 423680 3130 423732 3136
rect 424968 3188 425020 3194
rect 424968 3130 425020 3136
rect 424980 480 425008 3130
rect 428476 480 428504 11766
rect 432064 480 432092 15846
rect 442632 14476 442684 14482
rect 442632 14418 442684 14424
rect 439136 3324 439188 3330
rect 439136 3266 439188 3272
rect 435548 3256 435600 3262
rect 435548 3198 435600 3204
rect 435560 480 435588 3198
rect 439148 480 439176 3266
rect 442644 480 442672 14418
rect 552664 13116 552716 13122
rect 552664 13058 552716 13064
rect 470600 11756 470652 11762
rect 470600 11698 470652 11704
rect 449808 4140 449860 4146
rect 449808 4082 449860 4088
rect 446220 3392 446272 3398
rect 446220 3334 446272 3340
rect 446232 480 446260 3334
rect 449820 480 449848 4082
rect 453304 4072 453356 4078
rect 453304 4014 453356 4020
rect 453316 480 453344 4014
rect 456892 4004 456944 4010
rect 456892 3946 456944 3952
rect 456904 480 456932 3946
rect 460388 3936 460440 3942
rect 460388 3878 460440 3884
rect 460400 480 460428 3878
rect 467472 3868 467524 3874
rect 467472 3810 467524 3816
rect 463976 3800 464028 3806
rect 463976 3742 464028 3748
rect 463988 480 464016 3742
rect 467484 480 467512 3810
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 11698
rect 548616 10328 548668 10334
rect 548616 10270 548668 10276
rect 545488 8968 545540 8974
rect 545488 8910 545540 8916
rect 534906 7712 534962 7721
rect 527824 7676 527876 7682
rect 534906 7647 534962 7656
rect 527824 7618 527876 7624
rect 524236 6248 524288 6254
rect 524236 6190 524288 6196
rect 488816 5296 488868 5302
rect 488816 5238 488868 5244
rect 485226 3768 485282 3777
rect 481732 3732 481784 3738
rect 485226 3703 485282 3712
rect 481732 3674 481784 3680
rect 478144 3664 478196 3670
rect 478144 3606 478196 3612
rect 474556 3596 474608 3602
rect 474556 3538 474608 3544
rect 474568 480 474596 3538
rect 478156 480 478184 3606
rect 481744 480 481772 3674
rect 485240 480 485268 3703
rect 488828 480 488856 5238
rect 495900 5228 495952 5234
rect 495900 5170 495952 5176
rect 492312 3460 492364 3466
rect 492312 3402 492364 3408
rect 492324 480 492352 3402
rect 495912 480 495940 5170
rect 502984 5160 503036 5166
rect 502984 5102 503036 5108
rect 499394 3632 499450 3641
rect 499394 3567 499450 3576
rect 499408 480 499436 3567
rect 502996 480 503024 5102
rect 506480 5092 506532 5098
rect 506480 5034 506532 5040
rect 506492 480 506520 5034
rect 513564 5024 513616 5030
rect 513564 4966 513616 4972
rect 510068 3528 510120 3534
rect 510068 3470 510120 3476
rect 510080 480 510108 3470
rect 513576 480 513604 4966
rect 517150 3496 517206 3505
rect 517150 3431 517206 3440
rect 517164 480 517192 3431
rect 520738 3360 520794 3369
rect 520738 3295 520794 3304
rect 520752 480 520780 3295
rect 524248 480 524276 6190
rect 527836 480 527864 7618
rect 531320 7608 531372 7614
rect 531320 7550 531372 7556
rect 531332 480 531360 7550
rect 534920 480 534948 7647
rect 541990 7576 542046 7585
rect 541990 7511 542046 7520
rect 538404 6180 538456 6186
rect 538404 6122 538456 6128
rect 538416 480 538444 6122
rect 542004 480 542032 7511
rect 545500 480 545528 8910
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 10270
rect 552676 480 552704 13058
rect 556160 4956 556212 4962
rect 556160 4898 556212 4904
rect 556172 480 556200 4898
rect 559748 4888 559800 4894
rect 559748 4830 559800 4836
rect 559760 480 559788 4830
rect 562428 3466 562456 199378
rect 563244 4820 563296 4826
rect 563244 4762 563296 4768
rect 562416 3460 562468 3466
rect 562416 3402 562468 3408
rect 563256 480 563284 4762
rect 565096 3602 565124 242150
rect 565832 16574 565860 243510
rect 566476 126954 566504 453999
rect 569224 239420 569276 239426
rect 569224 239362 569276 239368
rect 566464 126948 566516 126954
rect 566464 126890 566516 126896
rect 565832 16546 566872 16574
rect 565084 3596 565136 3602
rect 565084 3538 565136 3544
rect 566844 480 566872 16546
rect 569236 3534 569264 239362
rect 569960 198008 570012 198014
rect 569960 197950 570012 197956
rect 569972 16574 570000 197950
rect 570616 167006 570644 454038
rect 570604 167000 570656 167006
rect 570604 166942 570656 166948
rect 571996 113150 572024 455495
rect 573376 153202 573404 455631
rect 580262 452704 580318 452713
rect 580262 452639 580318 452648
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 578884 236700 578936 236706
rect 578884 236642 578936 236648
rect 573364 153196 573416 153202
rect 573364 153138 573416 153144
rect 571984 113144 572036 113150
rect 571984 113086 572036 113092
rect 569972 16546 570368 16574
rect 569224 3528 569276 3534
rect 569224 3470 569276 3476
rect 570340 480 570368 16546
rect 573916 3596 573968 3602
rect 573916 3538 573968 3544
rect 573928 480 573956 3538
rect 577412 3528 577464 3534
rect 577412 3470 577464 3476
rect 577424 480 577452 3470
rect 578896 3126 578924 236642
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579988 113144 580040 113150
rect 579988 113086 580040 113092
rect 580000 112849 580028 113086
rect 579986 112840 580042 112849
rect 579986 112775 580042 112784
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580276 6633 580304 452639
rect 580368 99521 580396 458215
rect 580460 179217 580488 458254
rect 580446 179208 580502 179217
rect 580446 179143 580502 179152
rect 580552 139369 580580 458351
rect 580644 219065 580672 460906
rect 580724 458244 580776 458250
rect 580724 458186 580776 458192
rect 580736 232393 580764 458186
rect 580908 449540 580960 449546
rect 580908 449482 580960 449488
rect 580816 442264 580868 442270
rect 580816 442206 580868 442212
rect 580828 431633 580856 442206
rect 580814 431624 580870 431633
rect 580814 431559 580870 431568
rect 580816 422952 580868 422958
rect 580816 422894 580868 422900
rect 580828 298761 580856 422894
rect 580920 404977 580948 449482
rect 580906 404968 580962 404977
rect 580906 404903 580962 404912
rect 580814 298752 580870 298761
rect 580814 298687 580870 298696
rect 582380 247716 582432 247722
rect 582380 247658 582432 247664
rect 580722 232384 580778 232393
rect 580722 232319 580778 232328
rect 580630 219056 580686 219065
rect 580630 218991 580686 219000
rect 580814 194032 580870 194041
rect 580814 193967 580870 193976
rect 580630 193896 580686 193905
rect 580630 193831 580686 193840
rect 580538 139360 580594 139369
rect 580538 139295 580594 139304
rect 580446 105632 580502 105641
rect 580446 105567 580502 105576
rect 580354 99512 580410 99521
rect 580354 99447 580410 99456
rect 580460 59673 580488 105567
rect 580446 59664 580502 59673
rect 580446 59599 580502 59608
rect 580644 19825 580672 193831
rect 580722 105496 580778 105505
rect 580722 105431 580778 105440
rect 580736 73001 580764 105431
rect 580722 72992 580778 73001
rect 580722 72927 580778 72936
rect 580828 33153 580856 193967
rect 580906 105768 580962 105777
rect 580906 105703 580962 105712
rect 580920 86193 580948 105703
rect 580906 86184 580962 86193
rect 580906 86119 580962 86128
rect 580814 33144 580870 33153
rect 580814 33079 580870 33088
rect 580630 19816 580686 19825
rect 580630 19751 580686 19760
rect 582392 16574 582420 247658
rect 582392 16546 583432 16574
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 578884 3120 578936 3126
rect 578884 3062 578936 3068
rect 581000 3120 581052 3126
rect 581000 3062 581052 3068
rect 581012 480 581040 3062
rect 582208 480 582236 3402
rect 583404 480 583432 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 72974 700304 73030 700360
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658164 3478 658200
rect 3422 658144 3424 658164
rect 3424 658144 3476 658164
rect 3476 658144 3478 658164
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3330 501744 3386 501800
rect 3514 514800 3570 514856
rect 3054 475632 3110 475688
rect 3422 462576 3478 462632
rect 150990 674892 151046 674928
rect 150990 674872 150992 674892
rect 150992 674872 151044 674892
rect 151044 674872 151046 674892
rect 17590 626864 17646 626920
rect 17222 622784 17278 622840
rect 16026 587152 16082 587208
rect 3422 452240 3478 452296
rect 3330 449520 3386 449576
rect 3330 397432 3386 397488
rect 3054 371320 3110 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 2962 319232 3018 319288
rect 3330 306176 3386 306232
rect 2870 293120 2926 293176
rect 3238 267144 3294 267200
rect 3330 254088 3386 254144
rect 3238 241032 3294 241088
rect 3330 214920 3386 214976
rect 3330 201864 3386 201920
rect 3330 188808 3386 188864
rect 3054 136720 3110 136776
rect 3330 110608 3386 110664
rect 3330 71576 3386 71632
rect 3330 58520 3386 58576
rect 3330 45500 3332 45520
rect 3332 45500 3384 45520
rect 3384 45500 3386 45520
rect 3330 45464 3386 45500
rect 3330 32408 3386 32464
rect 3698 410488 3754 410544
rect 3606 162832 3662 162888
rect 3790 149776 3846 149832
rect 3698 84632 3754 84688
rect 14554 449928 14610 449984
rect 3514 19352 3570 19408
rect 15934 521464 15990 521520
rect 16302 508272 16358 508328
rect 15934 474000 15990 474056
rect 16946 533704 17002 533760
rect 17406 619928 17462 619984
rect 17314 599936 17370 599992
rect 17222 532752 17278 532808
rect 17498 618160 17554 618216
rect 17682 625912 17738 625968
rect 17590 536832 17646 536888
rect 17866 623736 17922 623792
rect 17774 621016 17830 621072
rect 17682 535880 17738 535936
rect 17590 532752 17646 532808
rect 17498 528128 17554 528184
rect 17498 527176 17554 527232
rect 16762 146920 16818 146976
rect 19246 598304 19302 598360
rect 19154 587696 19210 587752
rect 17866 533704 17922 533760
rect 17774 530984 17830 531040
rect 16946 144744 17002 144800
rect 16854 140800 16910 140856
rect 16670 139984 16726 140040
rect 17038 119992 17094 120048
rect 17314 146920 17370 146976
rect 17222 118360 17278 118416
rect 17038 29960 17094 30016
rect 17406 145968 17462 146024
rect 17314 56888 17370 56944
rect 17682 145968 17738 146024
rect 17682 144744 17738 144800
rect 17682 143792 17738 143848
rect 17590 142840 17646 142896
rect 17406 55936 17462 55992
rect 17590 139984 17646 140040
rect 17498 52808 17554 52864
rect 17774 140800 17830 140856
rect 17682 53760 17738 53816
rect 17866 138252 17868 138272
rect 17868 138252 17920 138272
rect 17920 138252 17922 138272
rect 17866 138216 17922 138252
rect 17774 51040 17830 51096
rect 17590 49952 17646 50008
rect 18786 529896 18842 529952
rect 36634 587832 36690 587888
rect 39578 587832 39634 587888
rect 42798 587832 42854 587888
rect 44178 587832 44234 587888
rect 45282 587832 45338 587888
rect 46846 587832 46902 587888
rect 48134 587832 48190 587888
rect 48686 587832 48742 587888
rect 49790 587832 49846 587888
rect 51078 587852 51134 587888
rect 51078 587832 51080 587852
rect 51080 587832 51132 587852
rect 51132 587832 51134 587852
rect 19338 536832 19394 536888
rect 19246 509904 19302 509960
rect 19154 491136 19210 491192
rect 18786 452784 18842 452840
rect 18602 449792 18658 449848
rect 18786 118088 18842 118144
rect 18418 107208 18474 107264
rect 17866 48184 17922 48240
rect 17222 28328 17278 28384
rect 18694 17312 18750 17368
rect 19430 508034 19486 508090
rect 48594 587696 48650 587752
rect 52366 587832 52422 587888
rect 53654 587832 53710 587888
rect 53838 587832 53894 587888
rect 55678 587832 55734 587888
rect 56230 587832 56286 587888
rect 59266 587832 59322 587888
rect 60554 587832 60610 587888
rect 61290 587832 61346 587888
rect 62762 587832 62818 587888
rect 63866 587832 63922 587888
rect 64970 587832 65026 587888
rect 66258 587832 66314 587888
rect 67638 587832 67694 587888
rect 68650 587832 68706 587888
rect 69754 587852 69810 587888
rect 69754 587832 69756 587852
rect 69756 587832 69808 587852
rect 69808 587832 69810 587852
rect 50066 587716 50122 587752
rect 50066 587696 50068 587716
rect 50068 587696 50120 587716
rect 50120 587696 50122 587716
rect 52642 587696 52698 587752
rect 57058 587424 57114 587480
rect 59818 587696 59874 587752
rect 61842 587288 61898 587344
rect 65522 587696 65578 587752
rect 65522 587424 65578 587480
rect 65982 587424 66038 587480
rect 63958 587288 64014 587344
rect 71134 587832 71190 587888
rect 72146 587832 72202 587888
rect 73250 587832 73306 587888
rect 73710 587832 73766 587888
rect 74354 587832 74410 587888
rect 76102 587832 76158 587888
rect 77390 587832 77446 587888
rect 78494 587832 78550 587888
rect 79138 587832 79194 587888
rect 81070 587832 81126 587888
rect 83646 587832 83702 587888
rect 88246 587832 88302 587888
rect 91006 587832 91062 587888
rect 93582 587832 93638 587888
rect 96066 587832 96122 587888
rect 98550 587832 98606 587888
rect 100942 587832 100998 587888
rect 103610 587832 103666 587888
rect 105542 587832 105598 587888
rect 108394 587832 108450 587888
rect 111246 587832 111302 587888
rect 113822 587832 113878 587888
rect 114558 587832 114614 587888
rect 118146 587832 118202 587888
rect 120538 587832 120594 587888
rect 125966 587832 126022 587888
rect 68558 587424 68614 587480
rect 122930 587016 122986 587072
rect 150714 585248 150770 585304
rect 122930 584568 122986 584624
rect 120538 584432 120594 584488
rect 118146 584296 118202 584352
rect 45374 499568 45430 499624
rect 37278 498072 37334 498128
rect 41878 498072 41934 498128
rect 43442 498072 43498 498128
rect 36174 497800 36230 497856
rect 37186 497820 37242 497856
rect 37186 497800 37188 497820
rect 37188 497800 37240 497820
rect 37240 497800 37242 497820
rect 22098 497564 22100 497584
rect 22100 497564 22152 497584
rect 22152 497564 22154 497584
rect 22098 497528 22154 497564
rect 19154 17448 19210 17504
rect 19798 107480 19854 107536
rect 18970 17176 19026 17232
rect 37278 491136 37334 491192
rect 39670 496984 39726 497040
rect 40590 496868 40646 496904
rect 40590 496848 40592 496868
rect 40592 496848 40644 496868
rect 40644 496848 40646 496868
rect 41878 494672 41934 494728
rect 44178 497936 44234 497992
rect 46846 498092 46902 498128
rect 46846 498072 46848 498092
rect 46848 498072 46900 498092
rect 46900 498072 46902 498092
rect 47582 498072 47638 498128
rect 48686 498072 48742 498128
rect 51446 498072 51502 498128
rect 52182 498108 52184 498128
rect 52184 498108 52236 498128
rect 52236 498108 52238 498128
rect 52182 498072 52238 498108
rect 53470 498072 53526 498128
rect 53838 498072 53894 498128
rect 55862 498072 55918 498128
rect 50250 497800 50306 497856
rect 57058 497800 57114 497856
rect 59542 498108 59544 498128
rect 59544 498108 59596 498128
rect 59596 498108 59598 498128
rect 59542 498072 59598 498108
rect 60646 498072 60702 498128
rect 63682 498072 63738 498128
rect 64142 498072 64198 498128
rect 67638 498072 67694 498128
rect 71226 498072 71282 498128
rect 71962 498072 72018 498128
rect 73710 498072 73766 498128
rect 73986 498072 74042 498128
rect 78126 498108 78128 498128
rect 78128 498108 78180 498128
rect 78180 498108 78182 498128
rect 78126 498072 78182 498108
rect 114466 498072 114522 498128
rect 121366 498072 121422 498128
rect 58162 497936 58218 497992
rect 61842 496984 61898 497040
rect 48318 496848 48374 496904
rect 50986 496848 51042 496904
rect 53746 496848 53802 496904
rect 56506 496848 56562 496904
rect 59266 496848 59322 496904
rect 62026 496848 62082 496904
rect 62762 496848 62818 496904
rect 68282 497120 68338 497176
rect 66258 496984 66314 497040
rect 65522 496868 65578 496904
rect 65522 496848 65524 496868
rect 65524 496848 65576 496868
rect 65576 496848 65578 496868
rect 66166 496848 66222 496904
rect 68558 496848 68614 496904
rect 73158 497700 73160 497720
rect 73160 497700 73212 497720
rect 73212 497700 73214 497720
rect 73158 497664 73214 497700
rect 69662 496848 69718 496904
rect 71686 496848 71742 496904
rect 76562 497936 76618 497992
rect 75182 497800 75238 497856
rect 73802 496848 73858 496904
rect 76838 496848 76894 496904
rect 78586 496848 78642 496904
rect 106094 497120 106150 497176
rect 79414 496848 79470 496904
rect 81346 496848 81402 496904
rect 84106 496848 84162 496904
rect 86866 496848 86922 496904
rect 88246 496848 88302 496904
rect 91006 496848 91062 496904
rect 93766 496848 93822 496904
rect 96526 496848 96582 496904
rect 99286 496848 99342 496904
rect 100942 496848 100998 496904
rect 104806 496848 104862 496904
rect 108854 496848 108910 496904
rect 111706 496848 111762 496904
rect 115846 496848 115902 496904
rect 118606 496848 118662 496904
rect 124126 496848 124182 496904
rect 126886 496848 126942 496904
rect 158718 668616 158774 668672
rect 157338 585656 157394 585712
rect 158718 579128 158774 579184
rect 156694 465704 156750 465760
rect 150990 196036 151046 196072
rect 150990 196016 150992 196036
rect 150992 196016 151044 196036
rect 151044 196016 151046 196036
rect 50802 109520 50858 109576
rect 56046 109520 56102 109576
rect 61106 109520 61162 109576
rect 106002 109520 106058 109576
rect 108578 109520 108634 109576
rect 48318 108976 48374 109032
rect 53654 108704 53710 108760
rect 68374 108976 68430 109032
rect 100942 108976 100998 109032
rect 111062 108976 111118 109032
rect 113454 108996 113510 109032
rect 113454 108976 113456 108996
rect 113456 108976 113508 108996
rect 113508 108976 113510 108996
rect 35898 107480 35954 107536
rect 36910 107516 36912 107536
rect 36912 107516 36964 107536
rect 36964 107516 36966 107536
rect 36910 107480 36966 107516
rect 38106 107480 38162 107536
rect 39578 107480 39634 107536
rect 40498 107480 40554 107536
rect 43166 107500 43222 107536
rect 43166 107480 43168 107500
rect 43168 107480 43220 107500
rect 43220 107480 43222 107500
rect 44270 107480 44326 107536
rect 45374 107480 45430 107536
rect 46570 107480 46626 107536
rect 47582 107480 47638 107536
rect 48778 107480 48834 107536
rect 50158 107516 50160 107536
rect 50160 107516 50212 107536
rect 50212 107516 50214 107536
rect 50158 107480 50214 107516
rect 51262 107480 51318 107536
rect 52366 107480 52422 107536
rect 53470 107480 53526 107536
rect 59634 107480 59690 107536
rect 60554 107480 60610 107536
rect 61658 107500 61714 107536
rect 61658 107480 61660 107500
rect 61660 107480 61712 107500
rect 61712 107480 61714 107500
rect 55126 107072 55182 107128
rect 55770 107072 55826 107128
rect 62578 107480 62634 107536
rect 63590 107480 63646 107536
rect 63866 107480 63922 107536
rect 65154 107480 65210 107536
rect 66258 107480 66314 107536
rect 67638 107480 67694 107536
rect 68650 107516 68652 107536
rect 68652 107516 68704 107536
rect 68704 107516 68706 107536
rect 68650 107480 68706 107516
rect 69754 107480 69810 107536
rect 71226 107480 71282 107536
rect 72146 107480 72202 107536
rect 73250 107480 73306 107536
rect 73710 107516 73712 107536
rect 73712 107516 73764 107536
rect 73764 107516 73766 107536
rect 73710 107480 73766 107516
rect 74354 107480 74410 107536
rect 75642 107500 75698 107536
rect 75642 107480 75644 107500
rect 75644 107480 75696 107500
rect 75696 107480 75698 107500
rect 61750 107344 61806 107400
rect 76102 107500 76158 107536
rect 76102 107480 76104 107500
rect 76104 107480 76156 107500
rect 76156 107480 76158 107500
rect 77666 107480 77722 107536
rect 78494 107480 78550 107536
rect 79138 107480 79194 107536
rect 86038 107480 86094 107536
rect 88246 107480 88302 107536
rect 93582 107480 93638 107536
rect 98550 107480 98606 107536
rect 120998 107480 121054 107536
rect 123390 107480 123446 107536
rect 57058 106256 57114 106312
rect 150806 105304 150862 105360
rect 52366 19488 52422 19544
rect 53470 19488 53526 19544
rect 55954 19488 56010 19544
rect 50894 18672 50950 18728
rect 36542 17892 36544 17912
rect 36544 17892 36596 17912
rect 36596 17892 36598 17912
rect 36542 17856 36598 17892
rect 43074 17856 43130 17912
rect 44178 17856 44234 17912
rect 45374 17856 45430 17912
rect 46662 17856 46718 17912
rect 47582 17856 47638 17912
rect 48686 17856 48742 17912
rect 50158 17856 50214 17912
rect 51446 17856 51502 17912
rect 19798 17584 19854 17640
rect 38658 17176 38714 17232
rect 53654 18692 53710 18728
rect 53654 18672 53656 18692
rect 53656 18672 53708 18692
rect 53708 18672 53710 18692
rect 95974 19216 96030 19272
rect 100942 19236 100998 19272
rect 100942 19216 100944 19236
rect 100944 19216 100996 19236
rect 100996 19216 100998 19236
rect 103702 19252 103704 19272
rect 103704 19252 103756 19272
rect 103756 19252 103758 19272
rect 103702 19216 103758 19252
rect 86038 19080 86094 19136
rect 91006 19100 91062 19136
rect 91006 19080 91008 19100
rect 91008 19080 91060 19100
rect 91060 19080 91062 19100
rect 76102 18944 76158 19000
rect 81070 18964 81126 19000
rect 81070 18944 81072 18964
rect 81072 18944 81124 18964
rect 81124 18944 81126 18964
rect 56046 18808 56102 18864
rect 58162 18828 58218 18864
rect 58162 18808 58164 18828
rect 58164 18808 58216 18828
rect 58216 18808 58218 18828
rect 73710 18828 73766 18864
rect 73710 18808 73712 18828
rect 73712 18808 73764 18828
rect 73764 18808 73766 18828
rect 106094 18556 106150 18592
rect 106094 18536 106096 18556
rect 106096 18536 106148 18556
rect 106148 18536 106150 18556
rect 108670 18536 108726 18592
rect 113454 18420 113510 18456
rect 113454 18400 113456 18420
rect 113456 18400 113508 18420
rect 113508 18400 113510 18420
rect 59542 17856 59598 17912
rect 60462 17876 60518 17912
rect 60462 17856 60464 17876
rect 60464 17856 60516 17876
rect 60516 17856 60518 17876
rect 53838 17584 53894 17640
rect 57886 17312 57942 17368
rect 62026 17892 62028 17912
rect 62028 17892 62080 17912
rect 62080 17892 62082 17912
rect 62026 17856 62082 17892
rect 64694 17876 64750 17912
rect 64694 17856 64696 17876
rect 64696 17856 64748 17876
rect 64748 17856 64750 17876
rect 66166 17856 66222 17912
rect 67638 17856 67694 17912
rect 71778 17856 71834 17912
rect 73158 17856 73214 17912
rect 78586 17856 78642 17912
rect 125966 17856 126022 17912
rect 68190 17584 68246 17640
rect 68926 17584 68982 17640
rect 70398 17584 70454 17640
rect 65062 17312 65118 17368
rect 66258 17332 66314 17368
rect 66258 17312 66260 17332
rect 66260 17312 66312 17332
rect 66312 17312 66314 17332
rect 69662 17448 69718 17504
rect 67638 17348 67640 17368
rect 67640 17348 67692 17368
rect 67692 17348 67694 17368
rect 67638 17312 67694 17348
rect 68190 17312 68246 17368
rect 60738 17176 60794 17232
rect 62118 17176 62174 17232
rect 63498 17196 63554 17232
rect 63498 17176 63500 17196
rect 63500 17176 63552 17196
rect 63552 17176 63554 17196
rect 69018 17176 69074 17232
rect 71686 17196 71742 17232
rect 71686 17176 71688 17196
rect 71688 17176 71740 17196
rect 71740 17176 71742 17196
rect 83830 17584 83886 17640
rect 75918 17448 75974 17504
rect 78678 17468 78734 17504
rect 78678 17448 78680 17468
rect 78680 17448 78732 17468
rect 78732 17448 78734 17468
rect 88246 17468 88302 17504
rect 88246 17448 88248 17468
rect 88248 17448 88300 17468
rect 88300 17448 88302 17468
rect 93582 17448 93638 17504
rect 99286 17332 99342 17368
rect 99286 17312 99288 17332
rect 99288 17312 99340 17332
rect 99340 17312 99342 17332
rect 111706 17312 111762 17368
rect 74814 17176 74870 17232
rect 77298 16924 77354 16960
rect 77298 16904 77300 16924
rect 77300 16904 77352 16924
rect 77352 16904 77354 16924
rect 173346 462984 173402 463040
rect 173162 462712 173218 462768
rect 170402 462576 170458 462632
rect 158718 189216 158774 189272
rect 158718 99184 158774 99240
rect 158902 99184 158958 99240
rect 173254 461216 173310 461272
rect 175922 462440 175978 462496
rect 173530 462304 173586 462360
rect 173530 19080 173586 19136
rect 173714 460944 173770 461000
rect 173806 456184 173862 456240
rect 173714 19216 173770 19272
rect 3422 6432 3478 6488
rect 176106 461080 176162 461136
rect 176014 459720 176070 459776
rect 179326 460264 179382 460320
rect 179142 459992 179198 460048
rect 178590 459856 178646 459912
rect 176198 459584 176254 459640
rect 176290 458632 176346 458688
rect 176474 458496 176530 458552
rect 176382 457544 176438 457600
rect 176566 452920 176622 452976
rect 178958 458768 179014 458824
rect 181810 457000 181866 457056
rect 182086 106664 182142 106720
rect 181442 17720 181498 17776
rect 184570 451560 184626 451616
rect 184662 450064 184718 450120
rect 185582 19080 185638 19136
rect 185490 18808 185546 18864
rect 186778 394712 186834 394768
rect 186318 247560 186374 247616
rect 187330 453328 187386 453384
rect 188342 451696 188398 451752
rect 188158 369008 188214 369064
rect 188342 18944 188398 19000
rect 188894 451424 188950 451480
rect 190090 451968 190146 452024
rect 189998 451832 190054 451888
rect 190826 398812 190882 398848
rect 190826 398792 190828 398812
rect 190828 398792 190880 398812
rect 190880 398792 190882 398812
rect 190826 397296 190882 397352
rect 190826 372564 190882 372600
rect 190826 372544 190828 372564
rect 190828 372544 190880 372564
rect 190880 372544 190882 372564
rect 191102 398792 191158 398848
rect 191102 397296 191158 397352
rect 188894 18672 188950 18728
rect 187422 17312 187478 17368
rect 195242 679360 195298 679416
rect 195334 679224 195390 679280
rect 195426 498072 195482 498128
rect 196438 678272 196494 678328
rect 196806 682080 196862 682136
rect 196990 679632 197046 679688
rect 196898 679088 196954 679144
rect 197818 465976 197874 466032
rect 191470 419600 191526 419656
rect 191470 397296 191526 397352
rect 191378 372544 191434 372600
rect 191378 369824 191434 369880
rect 198462 497664 198518 497720
rect 199290 679768 199346 679824
rect 199198 678136 199254 678192
rect 199474 679496 199530 679552
rect 201222 682216 201278 682272
rect 201130 681944 201186 682000
rect 197542 458360 197598 458416
rect 195978 458224 196034 458280
rect 196254 455504 196310 455560
rect 194598 454144 194654 454200
rect 193678 452648 193734 452704
rect 194506 450744 194562 450800
rect 194322 450472 194378 450528
rect 194506 450472 194562 450528
rect 194138 450200 194194 450256
rect 194322 450200 194378 450256
rect 195150 451424 195206 451480
rect 195886 451288 195942 451344
rect 197358 455640 197414 455696
rect 196990 454008 197046 454064
rect 201130 501608 201186 501664
rect 218978 700848 219034 700904
rect 201866 682760 201922 682816
rect 300122 700712 300178 700768
rect 332506 700576 332562 700632
rect 348790 700440 348846 700496
rect 364982 700304 365038 700360
rect 291106 682760 291162 682816
rect 238482 682624 238538 682680
rect 271970 682488 272026 682544
rect 274362 682352 274418 682408
rect 286322 682216 286378 682272
rect 283930 682080 283986 682136
rect 288714 681944 288770 682000
rect 305458 680448 305514 680504
rect 326986 682624 327042 682680
rect 319810 682488 319866 682544
rect 331770 680312 331826 680368
rect 341338 682216 341394 682272
rect 338946 682080 339002 682136
rect 367650 682352 367706 682408
rect 374826 682080 374882 682136
rect 372434 681944 372490 682000
rect 370042 681808 370098 681864
rect 209778 679768 209834 679824
rect 204994 679496 205050 679552
rect 264518 679632 264574 679688
rect 269302 679632 269358 679688
rect 300674 679496 300730 679552
rect 293498 679360 293554 679416
rect 295890 679224 295946 679280
rect 298282 679224 298338 679280
rect 212538 500248 212594 500304
rect 211158 500112 211214 500168
rect 201406 451424 201462 451480
rect 209870 480800 209926 480856
rect 211250 497392 211306 497448
rect 211342 462848 211398 462904
rect 211434 457408 211490 457464
rect 213918 500656 213974 500712
rect 214102 500656 214158 500712
rect 354862 500692 354864 500712
rect 354864 500692 354916 500712
rect 354916 500692 354918 500712
rect 212630 499840 212686 499896
rect 214010 500520 214066 500576
rect 215298 499976 215354 500032
rect 218058 468424 218114 468480
rect 228454 500384 228510 500440
rect 237654 498072 237710 498128
rect 234710 497528 234766 497584
rect 230110 453328 230166 453384
rect 232778 454280 232834 454336
rect 233422 449928 233478 449984
rect 234894 452240 234950 452296
rect 235998 452104 236054 452160
rect 320178 500520 320234 500576
rect 238942 497936 238998 497992
rect 288438 500384 288494 500440
rect 244922 499468 244924 499488
rect 244924 499468 244976 499488
rect 244976 499468 244978 499488
rect 244922 499432 244978 499468
rect 247038 497800 247094 497856
rect 245658 497664 245714 497720
rect 244462 494808 244518 494864
rect 245750 494672 245806 494728
rect 248602 466112 248658 466168
rect 248878 452512 248934 452568
rect 259734 494944 259790 495000
rect 277398 496032 277454 496088
rect 264702 451968 264758 452024
rect 265438 453192 265494 453248
rect 266174 451832 266230 451888
rect 266910 451696 266966 451752
rect 273258 463664 273314 463720
rect 272154 461352 272210 461408
rect 273902 453056 273958 453112
rect 280158 493312 280214 493368
rect 277674 454688 277730 454744
rect 283010 456864 283066 456920
rect 284206 451560 284262 451616
rect 284942 453056 284998 453112
rect 285954 457544 286010 457600
rect 230478 449792 230534 449848
rect 287702 474000 287758 474056
rect 287886 451288 287942 451344
rect 289082 454280 289138 454336
rect 290002 456184 290058 456240
rect 292302 451560 292358 451616
rect 298926 450608 298982 450664
rect 300398 452784 300454 452840
rect 300766 451832 300822 451888
rect 302330 462984 302386 463040
rect 304814 449928 304870 449984
rect 309322 458904 309378 458960
rect 310702 462712 310758 462768
rect 314658 465976 314714 466032
rect 314750 461216 314806 461272
rect 317418 465840 317474 465896
rect 316590 450472 316646 450528
rect 317510 462576 317566 462632
rect 319166 451696 319222 451752
rect 320638 450472 320694 450528
rect 329838 450336 329894 450392
rect 331402 460264 331458 460320
rect 332874 456048 332930 456104
rect 337658 459992 337714 460048
rect 338210 475360 338266 475416
rect 340510 450336 340566 450392
rect 342534 457272 342590 457328
rect 343914 459856 343970 459912
rect 354862 500656 354918 500692
rect 364154 500692 364156 500712
rect 364156 500692 364208 500712
rect 364208 500692 364210 500712
rect 346858 458768 346914 458824
rect 348330 455912 348386 455968
rect 350078 452920 350134 452976
rect 352746 459720 352802 459776
rect 352286 451968 352342 452024
rect 354494 450064 354550 450120
rect 355690 458632 355746 458688
rect 364154 500656 364210 500692
rect 366362 500656 366418 500712
rect 357438 450200 357494 450256
rect 359002 459584 359058 459640
rect 361670 458496 361726 458552
rect 364430 462440 364486 462496
rect 364062 452104 364118 452160
rect 369122 499976 369178 500032
rect 368754 452104 368810 452160
rect 378138 584704 378194 584760
rect 377862 584432 377918 584488
rect 377770 499976 377826 500032
rect 370134 461080 370190 461136
rect 369950 452376 370006 452432
rect 371882 457136 371938 457192
rect 373630 454552 373686 454608
rect 373262 452512 373318 452568
rect 372434 451832 372490 451888
rect 372434 450744 372490 450800
rect 372526 450608 372582 450664
rect 375102 455776 375158 455832
rect 375470 460944 375526 461000
rect 376206 452512 376262 452568
rect 375838 452240 375894 452296
rect 376850 461624 376906 461680
rect 377770 457000 377826 457056
rect 378138 451968 378194 452024
rect 378782 451832 378838 451888
rect 379058 584704 379114 584760
rect 379058 584568 379114 584624
rect 379610 462304 379666 462360
rect 379702 461488 379758 461544
rect 382554 460128 382610 460184
rect 382370 454416 382426 454472
rect 383658 450880 383714 450936
rect 389178 682080 389234 682136
rect 388166 681944 388222 682000
rect 385130 465704 385186 465760
rect 367006 449792 367062 449848
rect 261390 449656 261446 449712
rect 383934 449656 383990 449712
rect 387614 449520 387670 449576
rect 194046 449248 194102 449304
rect 191838 422320 191894 422376
rect 191838 419600 191894 419656
rect 191838 397296 191894 397352
rect 191838 395936 191894 395992
rect 191838 369144 191894 369200
rect 191838 369008 191894 369064
rect 191378 17448 191434 17504
rect 197358 247696 197414 247752
rect 201682 248240 201738 248296
rect 208398 247424 208454 247480
rect 213182 247832 213238 247888
rect 214562 247968 214618 248024
rect 215942 247288 215998 247344
rect 217322 249056 217378 249112
rect 216678 56888 216734 56944
rect 216678 55936 216734 55992
rect 216678 53780 216734 53816
rect 216678 53760 216680 53780
rect 216680 53760 216732 53780
rect 216732 53760 216734 53780
rect 216770 52808 216826 52864
rect 216770 51040 216826 51096
rect 216678 49952 216734 50008
rect 216678 48220 216680 48240
rect 216680 48220 216732 48240
rect 216732 48220 216734 48240
rect 216678 48184 216734 48220
rect 217138 3576 217194 3632
rect 217322 28464 217378 28520
rect 217322 28328 217378 28384
rect 217230 3440 217286 3496
rect 219162 3848 219218 3904
rect 218886 3304 218942 3360
rect 222842 248104 222898 248160
rect 222290 247832 222346 247888
rect 220910 247560 220966 247616
rect 219806 3712 219862 3768
rect 223670 247968 223726 248024
rect 223026 247832 223082 247888
rect 226430 248240 226486 248296
rect 225786 247968 225842 248024
rect 225050 247696 225106 247752
rect 225602 247696 225658 247752
rect 228362 247560 228418 247616
rect 227810 247288 227866 247344
rect 229190 247424 229246 247480
rect 254030 248104 254086 248160
rect 258170 247968 258226 248024
rect 256790 247832 256846 247888
rect 260930 247696 260986 247752
rect 265070 247560 265126 247616
rect 336738 111016 336794 111072
rect 340970 247560 341026 247616
rect 343730 247832 343786 247888
rect 345110 247696 345166 247752
rect 342258 111152 342314 111208
rect 347870 247968 347926 248024
rect 351182 106120 351238 106176
rect 353390 247288 353446 247344
rect 356794 247832 356850 247888
rect 356150 247152 356206 247208
rect 354770 247016 354826 247072
rect 285954 19488 286010 19544
rect 244278 19252 244280 19272
rect 244280 19252 244332 19272
rect 244332 19252 244334 19272
rect 244278 19216 244334 19252
rect 245290 19216 245346 19272
rect 246394 19236 246450 19272
rect 246394 19216 246396 19236
rect 246396 19216 246448 19236
rect 246448 19216 246450 19236
rect 248234 19100 248290 19136
rect 248234 19080 248236 19100
rect 248236 19080 248288 19100
rect 248288 19080 248290 19100
rect 250074 19080 250130 19136
rect 247498 18964 247554 19000
rect 247498 18944 247500 18964
rect 247500 18944 247552 18964
rect 247552 18944 247554 18964
rect 250626 18944 250682 19000
rect 252282 18828 252338 18864
rect 252282 18808 252284 18828
rect 252284 18808 252336 18828
rect 252336 18808 252338 18828
rect 253570 18808 253626 18864
rect 255962 18692 256018 18728
rect 255962 18672 255964 18692
rect 255964 18672 256016 18692
rect 256016 18672 256018 18692
rect 258354 18672 258410 18728
rect 235998 18536 236054 18592
rect 243082 18556 243138 18592
rect 243082 18536 243084 18556
rect 243084 18536 243136 18556
rect 243136 18536 243138 18556
rect 273258 17856 273314 17912
rect 277398 17876 277454 17912
rect 277398 17856 277400 17876
rect 277400 17856 277452 17876
rect 277452 17856 277454 17876
rect 280158 17892 280160 17912
rect 280160 17892 280212 17912
rect 280212 17892 280214 17912
rect 280158 17856 280214 17892
rect 263598 17720 263654 17776
rect 264978 17740 265034 17776
rect 264978 17720 264980 17740
rect 264980 17720 265032 17740
rect 265032 17720 265034 17740
rect 259550 17584 259606 17640
rect 260838 17584 260894 17640
rect 270498 17604 270554 17640
rect 270498 17584 270500 17604
rect 270500 17584 270552 17604
rect 270552 17584 270554 17604
rect 259458 17448 259514 17504
rect 255318 17312 255374 17368
rect 256698 17312 256754 17368
rect 258078 17332 258134 17368
rect 258078 17312 258080 17332
rect 258080 17312 258132 17332
rect 258132 17312 258134 17332
rect 282918 17176 282974 17232
rect 251178 17060 251234 17096
rect 251178 17040 251180 17060
rect 251180 17040 251232 17060
rect 251232 17040 251234 17060
rect 276018 3848 276074 3904
rect 279514 3712 279570 3768
rect 283102 3576 283158 3632
rect 286598 3440 286654 3496
rect 290186 3304 290242 3360
rect 357162 247288 357218 247344
rect 356978 247016 357034 247072
rect 358082 247968 358138 248024
rect 358266 247696 358322 247752
rect 358910 247016 358966 247072
rect 359738 99184 359794 99240
rect 360106 99184 360162 99240
rect 360842 247560 360898 247616
rect 388442 587152 388498 587208
rect 388442 450472 388498 450528
rect 388718 449928 388774 449984
rect 390558 681808 390614 681864
rect 388718 107344 388774 107400
rect 388534 106664 388590 106720
rect 388442 17720 388498 17776
rect 390374 451424 390430 451480
rect 391202 497392 391258 497448
rect 390190 142704 390246 142760
rect 390098 107072 390154 107128
rect 393962 462848 394018 462904
rect 407854 533296 407910 533352
rect 407762 500248 407818 500304
rect 399666 18808 399722 18864
rect 402334 19488 402390 19544
rect 402242 18672 402298 18728
rect 405002 17584 405058 17640
rect 405462 450336 405518 450392
rect 462318 700440 462374 700496
rect 543462 700304 543518 700360
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 551006 674892 551062 674928
rect 551006 674872 551008 674892
rect 551008 674872 551060 674892
rect 551060 674872 551062 674892
rect 417514 626864 417570 626920
rect 417146 625912 417202 625968
rect 416778 598032 416834 598088
rect 413282 584704 413338 584760
rect 410522 500112 410578 500168
rect 405370 19352 405426 19408
rect 405186 17448 405242 17504
rect 407670 109112 407726 109168
rect 407854 108976 407910 109032
rect 407762 17312 407818 17368
rect 408038 451560 408094 451616
rect 408314 450744 408370 450800
rect 408130 450608 408186 450664
rect 408314 109248 408370 109304
rect 408222 108840 408278 108896
rect 407946 17176 408002 17232
rect 410614 451288 410670 451344
rect 415858 527176 415914 527232
rect 416042 500384 416098 500440
rect 417422 599936 417478 599992
rect 417146 535880 417202 535936
rect 416686 493992 416742 494048
rect 414754 3440 414810 3496
rect 414938 3304 414994 3360
rect 416870 530984 416926 531040
rect 416962 529896 417018 529952
rect 416870 509924 416926 509960
rect 416870 509904 416872 509924
rect 416872 509904 416924 509924
rect 416924 509904 416926 509924
rect 418066 623736 418122 623792
rect 417974 621016 418030 621072
rect 417606 619928 417662 619984
rect 417514 536832 417570 536888
rect 417514 533724 417570 533760
rect 417514 533704 417516 533724
rect 417516 533704 417568 533724
rect 417568 533704 417570 533724
rect 417698 586880 417754 586936
rect 417422 509904 417478 509960
rect 417422 508000 417478 508056
rect 417790 508272 417846 508328
rect 417422 463664 417478 463720
rect 416778 146940 416834 146976
rect 416778 146920 416780 146940
rect 416780 146920 416832 146940
rect 416832 146920 416834 146940
rect 417330 146920 417386 146976
rect 417146 143792 417202 143848
rect 416778 141072 416834 141128
rect 416778 140020 416780 140040
rect 416780 140020 416832 140040
rect 416832 140020 416834 140040
rect 416778 139984 416834 140020
rect 417238 139984 417294 140040
rect 417146 119992 417202 120048
rect 416870 28328 416926 28384
rect 416778 28056 416834 28112
rect 417514 141072 417570 141128
rect 417422 118088 417478 118144
rect 417330 56888 417386 56944
rect 417238 49952 417294 50008
rect 419446 598306 419502 598362
rect 436282 587832 436338 587888
rect 438122 587832 438178 587888
rect 439594 587832 439650 587888
rect 441618 587832 441674 587888
rect 443090 587832 443146 587888
rect 444194 587832 444250 587888
rect 445666 587832 445722 587888
rect 446494 587832 446550 587888
rect 447322 587832 447378 587888
rect 448518 587832 448574 587888
rect 449898 587832 449954 587888
rect 450634 587832 450690 587888
rect 453578 587832 453634 587888
rect 454590 587832 454646 587888
rect 456062 587832 456118 587888
rect 456798 587832 456854 587888
rect 457258 587832 457314 587888
rect 471242 587832 471298 587888
rect 472162 587832 472218 587888
rect 419170 587560 419226 587616
rect 418710 587424 418766 587480
rect 418066 533704 418122 533760
rect 417974 530984 418030 531040
rect 418986 587288 419042 587344
rect 417790 118360 417846 118416
rect 417606 53760 417662 53816
rect 417514 51040 417570 51096
rect 417422 29960 417478 30016
rect 417790 28328 417846 28384
rect 418710 496712 418766 496768
rect 418066 107480 418122 107536
rect 418434 19080 418490 19136
rect 419170 500520 419226 500576
rect 436282 584840 436338 584896
rect 452382 587696 452438 587752
rect 453486 587696 453542 587752
rect 451370 586880 451426 586936
rect 456154 587696 456210 587752
rect 456798 586880 456854 586936
rect 458270 587696 458326 587752
rect 460662 587696 460718 587752
rect 460938 587696 460994 587752
rect 461582 587696 461638 587752
rect 462318 587696 462374 587752
rect 463882 587696 463938 587752
rect 465078 587696 465134 587752
rect 466274 587696 466330 587752
rect 467562 587696 467618 587752
rect 468666 587696 468722 587752
rect 469770 587696 469826 587752
rect 458178 587152 458234 587208
rect 462778 587188 462780 587208
rect 462780 587188 462832 587208
rect 462832 587188 462834 587208
rect 462778 587152 462834 587188
rect 460938 584704 460994 584760
rect 465170 587152 465226 587208
rect 473358 587832 473414 587888
rect 473634 587832 473690 587888
rect 476946 587852 477002 587888
rect 476946 587832 476948 587852
rect 476948 587832 477000 587852
rect 477000 587832 477002 587852
rect 473266 587696 473322 587752
rect 478050 587832 478106 587888
rect 479154 587832 479210 587888
rect 480258 587832 480314 587888
rect 483018 587832 483074 587888
rect 485778 587832 485834 587888
rect 487158 587832 487214 587888
rect 492678 587832 492734 587888
rect 495438 587832 495494 587888
rect 498198 587832 498254 587888
rect 500958 587832 501014 587888
rect 502338 587832 502394 587888
rect 505098 587832 505154 587888
rect 507858 587832 507914 587888
rect 510618 587832 510674 587888
rect 513378 587832 513434 587888
rect 514758 587832 514814 587888
rect 520278 587832 520334 587888
rect 470598 586472 470654 586528
rect 465078 584568 465134 584624
rect 489918 586472 489974 586528
rect 507858 584432 507914 584488
rect 523314 587832 523370 587888
rect 525890 587852 525946 587888
rect 525890 587832 525892 587852
rect 525892 587832 525944 587852
rect 525944 587832 525946 587852
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 558918 668616 558974 668672
rect 550822 585248 550878 585304
rect 514758 584296 514814 584352
rect 558918 579128 558974 579184
rect 441618 498072 441674 498128
rect 445298 498072 445354 498128
rect 449162 498072 449218 498128
rect 451278 498072 451334 498128
rect 452382 498072 452438 498128
rect 454590 498108 454592 498128
rect 454592 498108 454644 498128
rect 454644 498108 454646 498128
rect 454590 498072 454646 498108
rect 455510 498072 455566 498128
rect 469218 498072 469274 498128
rect 473358 498108 473360 498128
rect 473360 498108 473412 498128
rect 473412 498108 473414 498128
rect 473358 498072 473414 498108
rect 473542 498072 473598 498128
rect 480534 498072 480590 498128
rect 494702 498072 494758 498128
rect 504362 498072 504418 498128
rect 512642 498072 512698 498128
rect 519542 498072 519598 498128
rect 436190 497936 436246 497992
rect 436190 496984 436246 497040
rect 436098 496868 436154 496904
rect 436098 496848 436100 496868
rect 436100 496848 436152 496868
rect 436152 496848 436154 496868
rect 420734 496712 420790 496768
rect 418802 107208 418858 107264
rect 437478 496848 437534 496904
rect 438858 496848 438914 496904
rect 440238 496848 440294 496904
rect 444194 497392 444250 497448
rect 443642 496848 443698 496904
rect 441618 493992 441674 494048
rect 450542 497392 450598 497448
rect 446678 497120 446734 497176
rect 447782 496984 447838 497040
rect 447138 496848 447194 496904
rect 449898 496848 449954 496904
rect 453302 496984 453358 497040
rect 452658 496848 452714 496904
rect 463698 497936 463754 497992
rect 467838 497936 467894 497992
rect 460570 497800 460626 497856
rect 462318 497800 462374 497856
rect 457442 497392 457498 497448
rect 456062 496848 456118 496904
rect 456890 496848 456946 496904
rect 461122 497256 461178 497312
rect 462502 497392 462558 497448
rect 466458 497412 466514 497448
rect 466458 497392 466460 497412
rect 466460 497392 466512 497412
rect 466512 497392 466514 497412
rect 470874 497664 470930 497720
rect 465078 497276 465134 497312
rect 465078 497256 465080 497276
rect 465080 497256 465132 497276
rect 465132 497256 465134 497276
rect 465078 497120 465134 497176
rect 473358 497140 473414 497176
rect 473358 497120 473360 497140
rect 473360 497120 473412 497140
rect 473412 497120 473414 497140
rect 462042 496984 462098 497040
rect 471978 496984 472034 497040
rect 458178 496848 458234 496904
rect 459466 496868 459522 496904
rect 459466 496848 459468 496868
rect 459468 496848 459520 496868
rect 459520 496848 459522 496868
rect 460938 496848 460994 496904
rect 462410 496848 462466 496904
rect 465170 496848 465226 496904
rect 467930 496848 467986 496904
rect 470782 496848 470838 496904
rect 474738 497664 474794 497720
rect 476118 497684 476174 497720
rect 476118 497664 476120 497684
rect 476120 497664 476172 497684
rect 476172 497664 476174 497684
rect 478878 497256 478934 497312
rect 477590 496984 477646 497040
rect 476118 496848 476174 496904
rect 477498 496868 477554 496904
rect 477498 496848 477500 496868
rect 477500 496848 477552 496868
rect 477552 496848 477554 496868
rect 483018 496848 483074 496904
rect 485778 496848 485834 496904
rect 487158 496848 487214 496904
rect 490470 496848 490526 496904
rect 492678 496848 492734 496904
rect 497462 496848 497518 496904
rect 500958 496848 501014 496904
rect 502338 496848 502394 496904
rect 507858 496848 507914 496904
rect 510618 496848 510674 496904
rect 514758 496848 514814 496904
rect 517518 496848 517574 496904
rect 523038 496848 523094 496904
rect 525798 496848 525854 496904
rect 558182 454144 558238 454200
rect 551006 196036 551062 196072
rect 551006 196016 551008 196036
rect 551008 196016 551060 196036
rect 551060 196016 551062 196036
rect 451278 109792 451334 109848
rect 480902 109792 480958 109848
rect 483478 109792 483534 109848
rect 485962 109792 486018 109848
rect 488262 109792 488318 109848
rect 491022 109792 491078 109848
rect 436098 107480 436154 107536
rect 437018 107480 437074 107536
rect 438122 107480 438178 107536
rect 439594 107480 439650 107536
rect 440514 107480 440570 107536
rect 441618 107480 441674 107536
rect 443090 107480 443146 107536
rect 444194 107480 444250 107536
rect 445666 107480 445722 107536
rect 446402 107480 446458 107536
rect 447138 107480 447194 107536
rect 448518 107480 448574 107536
rect 449898 107480 449954 107536
rect 450634 107480 450690 107536
rect 476118 109656 476174 109712
rect 456982 109520 457038 109576
rect 493414 109656 493470 109712
rect 495898 109656 495954 109712
rect 498474 109656 498530 109712
rect 505926 109520 505982 109576
rect 508502 109520 508558 109576
rect 515862 109520 515918 109576
rect 518438 109520 518494 109576
rect 500958 108976 501014 109032
rect 503442 108976 503498 109032
rect 513378 108976 513434 109032
rect 457994 108432 458050 108488
rect 520922 108976 520978 109032
rect 523314 108976 523370 109032
rect 525890 108976 525946 109032
rect 452566 107480 452622 107536
rect 453578 107480 453634 107536
rect 454590 107480 454646 107536
rect 455786 107480 455842 107536
rect 455970 107500 456026 107536
rect 455970 107480 455972 107500
rect 455972 107480 456024 107500
rect 456024 107480 456026 107500
rect 453946 107072 454002 107128
rect 458362 107516 458364 107536
rect 458364 107516 458416 107536
rect 458416 107516 458418 107536
rect 458362 107480 458418 107516
rect 459466 107480 459522 107536
rect 460662 107480 460718 107536
rect 461674 107480 461730 107536
rect 462778 107480 462834 107536
rect 463882 107480 463938 107536
rect 465170 107480 465226 107536
rect 465722 107480 465778 107536
rect 467010 107480 467066 107536
rect 468666 107480 468722 107536
rect 469770 107480 469826 107536
rect 471150 107480 471206 107536
rect 472070 107480 472126 107536
rect 473358 107480 473414 107536
rect 474370 107500 474426 107536
rect 474370 107480 474372 107500
rect 474372 107480 474424 107500
rect 474424 107480 474426 107500
rect 457994 107072 458050 107128
rect 475658 107480 475714 107536
rect 478050 107516 478052 107536
rect 478052 107516 478104 107536
rect 478104 107516 478106 107536
rect 478050 107480 478106 107516
rect 479154 107480 479210 107536
rect 550730 105304 550786 105360
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580538 458360 580594 458416
rect 580354 458224 580410 458280
rect 580170 458088 580226 458144
rect 573362 455640 573418 455696
rect 571982 455504 572038 455560
rect 566462 454008 566518 454064
rect 558918 189080 558974 189136
rect 558918 99320 558974 99376
rect 460662 19780 460718 19816
rect 460662 19760 460664 19780
rect 460664 19760 460716 19780
rect 460716 19760 460718 19780
rect 488262 19760 488318 19816
rect 447598 19624 447654 19680
rect 448702 19624 448758 19680
rect 450082 19624 450138 19680
rect 455970 19624 456026 19680
rect 436098 17856 436154 17912
rect 436282 17856 436338 17912
rect 437478 17856 437534 17912
rect 438858 17856 438914 17912
rect 440238 17856 440294 17912
rect 441710 17856 441766 17912
rect 443090 17856 443146 17912
rect 444286 17876 444342 17912
rect 444286 17856 444288 17876
rect 444288 17856 444340 17876
rect 444340 17856 444342 17876
rect 445666 17856 445722 17912
rect 446494 17856 446550 17912
rect 447138 17856 447194 17912
rect 449898 17856 449954 17912
rect 451278 17856 451334 17912
rect 452290 17856 452346 17912
rect 453486 17856 453542 17912
rect 454038 17856 454094 17912
rect 455418 17856 455474 17912
rect 458362 17992 458418 18048
rect 473358 19624 473414 19680
rect 468298 19488 468354 19544
rect 470874 18808 470930 18864
rect 457350 17856 457406 17912
rect 458086 17856 458142 17912
rect 458270 17856 458326 17912
rect 459466 17856 459522 17912
rect 462318 17876 462374 17912
rect 462318 17856 462320 17876
rect 462320 17856 462372 17876
rect 462372 17856 462374 17876
rect 463698 17856 463754 17912
rect 465078 17856 465134 17912
rect 466458 17856 466514 17912
rect 467838 17856 467894 17912
rect 473358 17856 473414 17912
rect 471702 17312 471758 17368
rect 471978 17176 472034 17232
rect 465078 17040 465134 17096
rect 469310 17040 469366 17096
rect 471702 17040 471758 17096
rect 470874 16788 470930 16824
rect 470874 16768 470876 16788
rect 470876 16768 470928 16788
rect 470928 16768 470930 16788
rect 491022 19644 491078 19680
rect 491022 19624 491024 19644
rect 491024 19624 491076 19644
rect 491076 19624 491078 19644
rect 493414 19624 493470 19680
rect 495898 19508 495954 19544
rect 495898 19488 495900 19508
rect 495900 19488 495952 19508
rect 495952 19488 495954 19508
rect 500958 19488 501014 19544
rect 503534 19488 503590 19544
rect 485042 19216 485098 19272
rect 498474 19216 498530 19272
rect 501050 19216 501106 19272
rect 485042 18808 485098 18864
rect 515770 18964 515826 19000
rect 515770 18944 515772 18964
rect 515772 18944 515824 18964
rect 515824 18944 515826 18964
rect 501050 18808 501106 18864
rect 505834 18844 505836 18864
rect 505836 18844 505888 18864
rect 505888 18844 505890 18864
rect 505834 18808 505890 18844
rect 508410 18828 508466 18864
rect 508410 18808 508412 18828
rect 508412 18808 508464 18828
rect 508464 18808 508466 18828
rect 523314 18692 523370 18728
rect 523314 18672 523316 18692
rect 523316 18672 523368 18692
rect 523368 18672 523370 18692
rect 525890 18672 525946 18728
rect 476118 17856 476174 17912
rect 478878 17892 478880 17912
rect 478880 17892 478932 17912
rect 478932 17892 478934 17912
rect 478878 17856 478934 17892
rect 475382 17720 475438 17776
rect 475382 17448 475438 17504
rect 474738 17176 474794 17232
rect 477498 16904 477554 16960
rect 534906 7656 534962 7712
rect 485226 3712 485282 3768
rect 499394 3576 499450 3632
rect 517150 3440 517206 3496
rect 520738 3304 520794 3360
rect 541990 7520 542046 7576
rect 580262 452648 580318 452704
rect 580170 418240 580226 418296
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 272176 580226 272232
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579802 205672 579858 205728
rect 579618 192480 579674 192536
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 125976 580226 126032
rect 579986 112784 580042 112840
rect 580170 46280 580226 46336
rect 580446 179152 580502 179208
rect 580814 431568 580870 431624
rect 580906 404912 580962 404968
rect 580814 298696 580870 298752
rect 580722 232328 580778 232384
rect 580630 219000 580686 219056
rect 580814 193976 580870 194032
rect 580630 193840 580686 193896
rect 580538 139304 580594 139360
rect 580446 105576 580502 105632
rect 580354 99456 580410 99512
rect 580446 59608 580502 59664
rect 580722 105440 580778 105496
rect 580722 72936 580778 72992
rect 580906 105712 580962 105768
rect 580906 86128 580962 86184
rect 580814 33088 580870 33144
rect 580630 19760 580686 19816
rect 580262 6568 580318 6624
<< metal3 >>
rect 203190 700844 203196 700908
rect 203260 700906 203266 700908
rect 218973 700906 219039 700909
rect 203260 700904 219039 700906
rect 203260 700848 218978 700904
rect 219034 700848 219039 700904
rect 203260 700846 219039 700848
rect 203260 700844 203266 700846
rect 218973 700843 219039 700846
rect 202454 700708 202460 700772
rect 202524 700770 202530 700772
rect 300117 700770 300183 700773
rect 202524 700768 300183 700770
rect 202524 700712 300122 700768
rect 300178 700712 300183 700768
rect 202524 700710 300183 700712
rect 202524 700708 202530 700710
rect 300117 700707 300183 700710
rect 202270 700572 202276 700636
rect 202340 700634 202346 700636
rect 332501 700634 332567 700637
rect 202340 700632 332567 700634
rect 202340 700576 332506 700632
rect 332562 700576 332567 700632
rect 202340 700574 332567 700576
rect 202340 700572 202346 700574
rect 332501 700571 332567 700574
rect 202086 700436 202092 700500
rect 202156 700498 202162 700500
rect 348785 700498 348851 700501
rect 202156 700496 348851 700498
rect 202156 700440 348790 700496
rect 348846 700440 348851 700496
rect 202156 700438 348851 700440
rect 202156 700436 202162 700438
rect 348785 700435 348851 700438
rect 415894 700436 415900 700500
rect 415964 700498 415970 700500
rect 462313 700498 462379 700501
rect 415964 700496 462379 700498
rect 415964 700440 462318 700496
rect 462374 700440 462379 700496
rect 415964 700438 462379 700440
rect 415964 700436 415970 700438
rect 462313 700435 462379 700438
rect 72969 700362 73035 700365
rect 199326 700362 199332 700364
rect 72969 700360 199332 700362
rect 72969 700304 72974 700360
rect 73030 700304 199332 700360
rect 72969 700302 199332 700304
rect 72969 700299 73035 700302
rect 199326 700300 199332 700302
rect 199396 700300 199402 700364
rect 202638 700300 202644 700364
rect 202708 700362 202714 700364
rect 364977 700362 365043 700365
rect 202708 700360 365043 700362
rect 202708 700304 364982 700360
rect 365038 700304 365043 700360
rect 202708 700302 365043 700304
rect 202708 700300 202714 700302
rect 364977 700299 365043 700302
rect 418654 700300 418660 700364
rect 418724 700362 418730 700364
rect 543457 700362 543523 700365
rect 418724 700360 543523 700362
rect 418724 700304 543462 700360
rect 543518 700304 543523 700360
rect 418724 700302 543523 700304
rect 418724 700300 418730 700302
rect 543457 700299 543523 700302
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 201861 682818 201927 682821
rect 291101 682818 291167 682821
rect 201861 682816 291167 682818
rect 201861 682760 201866 682816
rect 201922 682760 291106 682816
rect 291162 682760 291167 682816
rect 201861 682758 291167 682760
rect 201861 682755 201927 682758
rect 291101 682755 291167 682758
rect 203558 682620 203564 682684
rect 203628 682682 203634 682684
rect 238477 682682 238543 682685
rect 203628 682680 238543 682682
rect 203628 682624 238482 682680
rect 238538 682624 238543 682680
rect 203628 682622 238543 682624
rect 203628 682620 203634 682622
rect 238477 682619 238543 682622
rect 326981 682682 327047 682685
rect 374126 682682 374132 682684
rect 326981 682680 374132 682682
rect 326981 682624 326986 682680
rect 327042 682624 374132 682680
rect 326981 682622 374132 682624
rect 326981 682619 327047 682622
rect 374126 682620 374132 682622
rect 374196 682620 374202 682684
rect 203742 682484 203748 682548
rect 203812 682546 203818 682548
rect 271965 682546 272031 682549
rect 203812 682544 272031 682546
rect 203812 682488 271970 682544
rect 272026 682488 272031 682544
rect 203812 682486 272031 682488
rect 203812 682484 203818 682486
rect 271965 682483 272031 682486
rect 319805 682546 319871 682549
rect 375414 682546 375420 682548
rect 319805 682544 375420 682546
rect 319805 682488 319810 682544
rect 319866 682488 375420 682544
rect 319805 682486 375420 682488
rect 319805 682483 319871 682486
rect 375414 682484 375420 682486
rect 375484 682484 375490 682548
rect 203374 682348 203380 682412
rect 203444 682410 203450 682412
rect 274357 682410 274423 682413
rect 203444 682408 274423 682410
rect 203444 682352 274362 682408
rect 274418 682352 274423 682408
rect 203444 682350 274423 682352
rect 203444 682348 203450 682350
rect 274357 682347 274423 682350
rect 367645 682410 367711 682413
rect 378174 682410 378180 682412
rect 367645 682408 378180 682410
rect 367645 682352 367650 682408
rect 367706 682352 378180 682408
rect 367645 682350 378180 682352
rect 367645 682347 367711 682350
rect 378174 682348 378180 682350
rect 378244 682348 378250 682412
rect 201217 682274 201283 682277
rect 286317 682274 286383 682277
rect 201217 682272 286383 682274
rect 201217 682216 201222 682272
rect 201278 682216 286322 682272
rect 286378 682216 286383 682272
rect 201217 682214 286383 682216
rect 201217 682211 201283 682214
rect 286317 682211 286383 682214
rect 341333 682274 341399 682277
rect 373758 682274 373764 682276
rect 341333 682272 373764 682274
rect 341333 682216 341338 682272
rect 341394 682216 373764 682272
rect 341333 682214 373764 682216
rect 341333 682211 341399 682214
rect 373758 682212 373764 682214
rect 373828 682212 373834 682276
rect 196801 682138 196867 682141
rect 283925 682138 283991 682141
rect 196801 682136 283991 682138
rect 196801 682080 196806 682136
rect 196862 682080 283930 682136
rect 283986 682080 283991 682136
rect 196801 682078 283991 682080
rect 196801 682075 196867 682078
rect 283925 682075 283991 682078
rect 338941 682138 339007 682141
rect 372654 682138 372660 682140
rect 338941 682136 372660 682138
rect 338941 682080 338946 682136
rect 339002 682080 372660 682136
rect 338941 682078 372660 682080
rect 338941 682075 339007 682078
rect 372654 682076 372660 682078
rect 372724 682076 372730 682140
rect 374821 682138 374887 682141
rect 389173 682138 389239 682141
rect 374821 682136 389239 682138
rect 374821 682080 374826 682136
rect 374882 682080 389178 682136
rect 389234 682080 389239 682136
rect 374821 682078 389239 682080
rect 374821 682075 374887 682078
rect 389173 682075 389239 682078
rect 201125 682002 201191 682005
rect 288709 682002 288775 682005
rect 201125 682000 288775 682002
rect 201125 681944 201130 682000
rect 201186 681944 288714 682000
rect 288770 681944 288775 682000
rect 201125 681942 288775 681944
rect 201125 681939 201191 681942
rect 288709 681939 288775 681942
rect 372429 682002 372495 682005
rect 388161 682002 388227 682005
rect 372429 682000 388227 682002
rect 372429 681944 372434 682000
rect 372490 681944 388166 682000
rect 388222 681944 388227 682000
rect 372429 681942 388227 681944
rect 372429 681939 372495 681942
rect 388161 681939 388227 681942
rect 370037 681866 370103 681869
rect 390553 681866 390619 681869
rect 370037 681864 390619 681866
rect 370037 681808 370042 681864
rect 370098 681808 390558 681864
rect 390614 681808 390619 681864
rect 370037 681806 390619 681808
rect 370037 681803 370103 681806
rect 390553 681803 390619 681806
rect 199878 680444 199884 680508
rect 199948 680506 199954 680508
rect 305453 680506 305519 680509
rect 199948 680504 305519 680506
rect 199948 680448 305458 680504
rect 305514 680448 305519 680504
rect 199948 680446 305519 680448
rect 199948 680444 199954 680446
rect 305453 680443 305519 680446
rect 195830 680308 195836 680372
rect 195900 680370 195906 680372
rect 331765 680370 331831 680373
rect 195900 680368 331831 680370
rect 195900 680312 331770 680368
rect 331826 680312 331831 680368
rect 195900 680310 331831 680312
rect 195900 680308 195906 680310
rect 331765 680307 331831 680310
rect 199285 679826 199351 679829
rect 209773 679826 209839 679829
rect 199285 679824 209839 679826
rect 199285 679768 199290 679824
rect 199346 679768 209778 679824
rect 209834 679768 209839 679824
rect 199285 679766 209839 679768
rect 199285 679763 199351 679766
rect 209773 679763 209839 679766
rect 196985 679690 197051 679693
rect 264513 679692 264579 679693
rect 269297 679692 269363 679693
rect 264462 679690 264468 679692
rect 196985 679688 205650 679690
rect 196985 679632 196990 679688
rect 197046 679632 205650 679688
rect 196985 679630 205650 679632
rect 264422 679630 264468 679690
rect 264532 679688 264579 679692
rect 269246 679690 269252 679692
rect 264574 679632 264579 679688
rect 196985 679627 197051 679630
rect 199469 679554 199535 679557
rect 204989 679554 205055 679557
rect 199469 679552 205055 679554
rect 199469 679496 199474 679552
rect 199530 679496 204994 679552
rect 205050 679496 205055 679552
rect 199469 679494 205055 679496
rect 205590 679554 205650 679630
rect 264462 679628 264468 679630
rect 264532 679628 264579 679632
rect 269206 679630 269252 679690
rect 269316 679688 269363 679692
rect 269358 679632 269363 679688
rect 269246 679628 269252 679630
rect 269316 679628 269363 679632
rect 264513 679627 264579 679628
rect 269297 679627 269363 679628
rect 300669 679554 300735 679557
rect 205590 679552 300735 679554
rect 205590 679496 300674 679552
rect 300730 679496 300735 679552
rect 205590 679494 300735 679496
rect 199469 679491 199535 679494
rect 204989 679491 205055 679494
rect 300669 679491 300735 679494
rect 195237 679418 195303 679421
rect 293493 679418 293559 679421
rect 195237 679416 293559 679418
rect 195237 679360 195242 679416
rect 195298 679360 293498 679416
rect 293554 679360 293559 679416
rect 195237 679358 293559 679360
rect 195237 679355 195303 679358
rect 293493 679355 293559 679358
rect 195329 679282 195395 679285
rect 295885 679282 295951 679285
rect 298277 679282 298343 679285
rect 195329 679280 295951 679282
rect 195329 679224 195334 679280
rect 195390 679224 295890 679280
rect 295946 679224 295951 679280
rect 195329 679222 295951 679224
rect 195329 679219 195395 679222
rect 295885 679219 295951 679222
rect 296670 679280 298343 679282
rect 296670 679224 298282 679280
rect 298338 679224 298343 679280
rect 296670 679222 298343 679224
rect 196893 679146 196959 679149
rect 296670 679146 296730 679222
rect 298277 679219 298343 679222
rect 196893 679144 296730 679146
rect 196893 679088 196898 679144
rect 196954 679088 296730 679144
rect 196893 679086 296730 679088
rect 196893 679083 196959 679086
rect 196433 678330 196499 678333
rect 264462 678330 264468 678332
rect 196433 678328 264468 678330
rect 196433 678272 196438 678328
rect 196494 678272 264468 678328
rect 196433 678270 264468 678272
rect 196433 678267 196499 678270
rect 264462 678268 264468 678270
rect 264532 678268 264538 678332
rect 199193 678194 199259 678197
rect 269246 678194 269252 678196
rect 199193 678192 269252 678194
rect 199193 678136 199198 678192
rect 199254 678136 269252 678192
rect 199193 678134 269252 678136
rect 199193 678131 199259 678134
rect 269246 678132 269252 678134
rect 269316 678132 269322 678196
rect 150985 674932 151051 674933
rect 551001 674932 551067 674933
rect 150934 674930 150940 674932
rect 150894 674870 150940 674930
rect 151004 674928 151051 674932
rect 550950 674930 550956 674932
rect 151046 674872 151051 674928
rect 150934 674868 150940 674870
rect 151004 674868 151051 674872
rect 550910 674870 550956 674930
rect 551020 674928 551067 674932
rect 551062 674872 551067 674928
rect 550950 674868 550956 674870
rect 551020 674868 551067 674872
rect 150985 674867 151051 674868
rect 551001 674867 551067 674868
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 156558 668674 156618 669190
rect 158713 668674 158779 668677
rect 156558 668672 158779 668674
rect 156558 668616 158718 668672
rect 158774 668616 158779 668672
rect 156558 668614 158779 668616
rect 556570 668674 556630 669190
rect 558913 668674 558979 668677
rect 556570 668672 558979 668674
rect 556570 668616 558918 668672
rect 558974 668616 558979 668672
rect 556570 668614 558979 668616
rect 158713 668611 158779 668614
rect 558913 668611 558979 668614
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 17585 626922 17651 626925
rect 19382 626922 20056 626924
rect 17585 626920 20056 626922
rect 17585 626864 17590 626920
rect 17646 626864 20056 626920
rect 417509 626922 417575 626925
rect 419398 626922 420072 626924
rect 417509 626920 420072 626922
rect 417509 626864 417514 626920
rect 417570 626864 420072 626920
rect 17585 626862 19442 626864
rect 417509 626862 419458 626864
rect 17585 626859 17651 626862
rect 417509 626859 417575 626862
rect 17677 625970 17743 625973
rect 19382 625970 20056 625972
rect 17677 625968 20056 625970
rect 17677 625912 17682 625968
rect 17738 625912 20056 625968
rect 417141 625970 417207 625973
rect 419398 625970 420072 625972
rect 417141 625968 420072 625970
rect 417141 625912 417146 625968
rect 417202 625912 420072 625968
rect 17677 625910 19442 625912
rect 417141 625910 419458 625912
rect 17677 625907 17743 625910
rect 417141 625907 417207 625910
rect 17861 623794 17927 623797
rect 19382 623794 20056 623796
rect 17861 623792 20056 623794
rect 17861 623736 17866 623792
rect 17922 623736 20056 623792
rect 418061 623794 418127 623797
rect 419398 623794 420072 623796
rect 418061 623792 420072 623794
rect 418061 623736 418066 623792
rect 418122 623736 420072 623792
rect 17861 623734 19442 623736
rect 418061 623734 419458 623736
rect 17861 623731 17927 623734
rect 418061 623731 418127 623734
rect 17217 622842 17283 622845
rect 19382 622842 20056 622844
rect 17217 622840 20056 622842
rect 17217 622784 17222 622840
rect 17278 622784 20056 622840
rect 17217 622782 19442 622784
rect 17217 622779 17283 622782
rect 417918 622780 417924 622844
rect 417988 622842 417994 622844
rect 419398 622842 420072 622844
rect 417988 622784 420072 622842
rect 417988 622782 419458 622784
rect 417988 622780 417994 622782
rect 17769 621074 17835 621077
rect 19382 621074 20056 621076
rect 17769 621072 20056 621074
rect 17769 621016 17774 621072
rect 17830 621016 20056 621072
rect 417969 621074 418035 621077
rect 419398 621074 420072 621076
rect 417969 621072 420072 621074
rect 417969 621016 417974 621072
rect 418030 621016 420072 621072
rect 17769 621014 19442 621016
rect 417969 621014 419458 621016
rect 17769 621011 17835 621014
rect 417969 621011 418035 621014
rect 17401 619986 17467 619989
rect 19382 619986 20056 619988
rect 17401 619984 20056 619986
rect 17401 619928 17406 619984
rect 17462 619928 20056 619984
rect 417601 619986 417667 619989
rect 419398 619986 420072 619988
rect 417601 619984 420072 619986
rect 417601 619928 417606 619984
rect 417662 619928 420072 619984
rect 17401 619926 19442 619928
rect 417601 619926 419458 619928
rect 17401 619923 17467 619926
rect 417601 619923 417667 619926
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 17493 618218 17559 618221
rect 19382 618218 20056 618220
rect 17493 618216 20056 618218
rect 17493 618160 17498 618216
rect 17554 618160 20056 618216
rect 17493 618158 19442 618160
rect 17493 618155 17559 618158
rect 417550 618156 417556 618220
rect 417620 618218 417626 618220
rect 419766 618218 420072 618220
rect 417620 618160 420072 618218
rect 417620 618158 419826 618160
rect 417620 618156 417626 618158
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect 17309 599994 17375 599997
rect 19382 599994 20056 599996
rect 17309 599992 20056 599994
rect 17309 599936 17314 599992
rect 17370 599936 20056 599992
rect 417417 599994 417483 599997
rect 419398 599994 420072 599996
rect 417417 599992 420072 599994
rect 417417 599936 417422 599992
rect 417478 599936 420072 599992
rect 17309 599934 19442 599936
rect 417417 599934 419458 599936
rect 17309 599931 17375 599934
rect 417417 599931 417483 599934
rect 19241 598362 19307 598365
rect 419441 598364 419507 598367
rect 19750 598362 20056 598364
rect 19241 598360 20056 598362
rect 19241 598304 19246 598360
rect 19302 598304 20056 598360
rect 419441 598362 420072 598364
rect 419441 598306 419446 598362
rect 419502 598306 420072 598362
rect 419441 598304 420072 598306
rect 19241 598302 19810 598304
rect 19241 598299 19307 598302
rect 419441 598301 419507 598304
rect 18638 598028 18644 598092
rect 18708 598090 18714 598092
rect 19382 598090 20056 598092
rect 18708 598032 20056 598090
rect 416773 598090 416839 598093
rect 419398 598090 420072 598092
rect 416773 598088 420072 598090
rect 416773 598032 416778 598088
rect 416834 598032 420072 598088
rect 18708 598030 19442 598032
rect 416773 598030 419458 598032
rect 18708 598028 18714 598030
rect 416773 598027 416839 598030
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 36629 587890 36695 587893
rect 39573 587892 39639 587893
rect 37038 587890 37044 587892
rect 36629 587888 37044 587890
rect 36629 587832 36634 587888
rect 36690 587832 37044 587888
rect 36629 587830 37044 587832
rect 36629 587827 36695 587830
rect 37038 587828 37044 587830
rect 37108 587828 37114 587892
rect 39573 587888 39620 587892
rect 39684 587890 39690 587892
rect 42793 587890 42859 587893
rect 44173 587892 44239 587893
rect 45277 587892 45343 587893
rect 43110 587890 43116 587892
rect 39573 587832 39578 587888
rect 39573 587828 39620 587832
rect 39684 587830 39730 587890
rect 42793 587888 43116 587890
rect 42793 587832 42798 587888
rect 42854 587832 43116 587888
rect 42793 587830 43116 587832
rect 39684 587828 39690 587830
rect 39573 587827 39639 587828
rect 42793 587827 42859 587830
rect 43110 587828 43116 587830
rect 43180 587828 43186 587892
rect 44173 587888 44220 587892
rect 44284 587890 44290 587892
rect 44173 587832 44178 587888
rect 44173 587828 44220 587832
rect 44284 587830 44330 587890
rect 45277 587888 45324 587892
rect 45388 587890 45394 587892
rect 45277 587832 45282 587888
rect 44284 587828 44290 587830
rect 45277 587828 45324 587832
rect 45388 587830 45434 587890
rect 45388 587828 45394 587830
rect 46606 587828 46612 587892
rect 46676 587890 46682 587892
rect 46841 587890 46907 587893
rect 46676 587888 46907 587890
rect 46676 587832 46846 587888
rect 46902 587832 46907 587888
rect 46676 587830 46907 587832
rect 46676 587828 46682 587830
rect 44173 587827 44239 587828
rect 45277 587827 45343 587828
rect 46841 587827 46907 587830
rect 47710 587828 47716 587892
rect 47780 587890 47786 587892
rect 48129 587890 48195 587893
rect 47780 587888 48195 587890
rect 47780 587832 48134 587888
rect 48190 587832 48195 587888
rect 47780 587830 48195 587832
rect 47780 587828 47786 587830
rect 48129 587827 48195 587830
rect 48262 587828 48268 587892
rect 48332 587890 48338 587892
rect 48681 587890 48747 587893
rect 48332 587888 48747 587890
rect 48332 587832 48686 587888
rect 48742 587832 48747 587888
rect 48332 587830 48747 587832
rect 48332 587828 48338 587830
rect 48681 587827 48747 587830
rect 49785 587890 49851 587893
rect 50654 587890 50660 587892
rect 49785 587888 50660 587890
rect 49785 587832 49790 587888
rect 49846 587832 50660 587888
rect 49785 587830 50660 587832
rect 49785 587827 49851 587830
rect 50654 587828 50660 587830
rect 50724 587828 50730 587892
rect 51073 587890 51139 587893
rect 52361 587892 52427 587893
rect 53649 587892 53715 587893
rect 51206 587890 51212 587892
rect 51073 587888 51212 587890
rect 51073 587832 51078 587888
rect 51134 587832 51212 587888
rect 51073 587830 51212 587832
rect 51073 587827 51139 587830
rect 51206 587828 51212 587830
rect 51276 587828 51282 587892
rect 52310 587890 52316 587892
rect 52270 587830 52316 587890
rect 52380 587888 52427 587892
rect 53598 587890 53604 587892
rect 52422 587832 52427 587888
rect 52310 587828 52316 587830
rect 52380 587828 52427 587832
rect 53558 587830 53604 587890
rect 53668 587888 53715 587892
rect 53710 587832 53715 587888
rect 53598 587828 53604 587830
rect 53668 587828 53715 587832
rect 52361 587827 52427 587828
rect 53649 587827 53715 587828
rect 53833 587890 53899 587893
rect 54518 587890 54524 587892
rect 53833 587888 54524 587890
rect 53833 587832 53838 587888
rect 53894 587832 54524 587888
rect 53833 587830 54524 587832
rect 53833 587827 53899 587830
rect 54518 587828 54524 587830
rect 54588 587828 54594 587892
rect 55673 587890 55739 587893
rect 55806 587890 55812 587892
rect 55673 587888 55812 587890
rect 55673 587832 55678 587888
rect 55734 587832 55812 587888
rect 55673 587830 55812 587832
rect 55673 587827 55739 587830
rect 55806 587828 55812 587830
rect 55876 587828 55882 587892
rect 55990 587828 55996 587892
rect 56060 587890 56066 587892
rect 56225 587890 56291 587893
rect 56060 587888 56291 587890
rect 56060 587832 56230 587888
rect 56286 587832 56291 587888
rect 56060 587830 56291 587832
rect 56060 587828 56066 587830
rect 56225 587827 56291 587830
rect 58566 587828 58572 587892
rect 58636 587890 58642 587892
rect 59261 587890 59327 587893
rect 58636 587888 59327 587890
rect 58636 587832 59266 587888
rect 59322 587832 59327 587888
rect 58636 587830 59327 587832
rect 58636 587828 58642 587830
rect 59261 587827 59327 587830
rect 60549 587892 60615 587893
rect 60549 587888 60596 587892
rect 60660 587890 60666 587892
rect 61285 587890 61351 587893
rect 62757 587892 62823 587893
rect 63861 587892 63927 587893
rect 61694 587890 61700 587892
rect 60549 587832 60554 587888
rect 60549 587828 60596 587832
rect 60660 587830 60706 587890
rect 61285 587888 61700 587890
rect 61285 587832 61290 587888
rect 61346 587832 61700 587888
rect 61285 587830 61700 587832
rect 60660 587828 60666 587830
rect 60549 587827 60615 587828
rect 61285 587827 61351 587830
rect 61694 587828 61700 587830
rect 61764 587828 61770 587892
rect 62757 587888 62804 587892
rect 62868 587890 62874 587892
rect 62757 587832 62762 587888
rect 62757 587828 62804 587832
rect 62868 587830 62914 587890
rect 63861 587888 63908 587892
rect 63972 587890 63978 587892
rect 64965 587890 65031 587893
rect 66253 587892 66319 587893
rect 67633 587892 67699 587893
rect 65190 587890 65196 587892
rect 63861 587832 63866 587888
rect 62868 587828 62874 587830
rect 63861 587828 63908 587832
rect 63972 587830 64018 587890
rect 64965 587888 65196 587890
rect 64965 587832 64970 587888
rect 65026 587832 65196 587888
rect 64965 587830 65196 587832
rect 63972 587828 63978 587830
rect 62757 587827 62823 587828
rect 63861 587827 63927 587828
rect 64965 587827 65031 587830
rect 65190 587828 65196 587830
rect 65260 587828 65266 587892
rect 66253 587888 66300 587892
rect 66364 587890 66370 587892
rect 67582 587890 67588 587892
rect 66253 587832 66258 587888
rect 66253 587828 66300 587832
rect 66364 587830 66410 587890
rect 67542 587830 67588 587890
rect 67652 587888 67699 587892
rect 67694 587832 67699 587888
rect 66364 587828 66370 587830
rect 67582 587828 67588 587830
rect 67652 587828 67699 587832
rect 66253 587827 66319 587828
rect 67633 587827 67699 587828
rect 68645 587892 68711 587893
rect 69749 587892 69815 587893
rect 68645 587888 68692 587892
rect 68756 587890 68762 587892
rect 68645 587832 68650 587888
rect 68645 587828 68692 587832
rect 68756 587830 68802 587890
rect 69749 587888 69796 587892
rect 69860 587890 69866 587892
rect 71129 587890 71195 587893
rect 72141 587892 72207 587893
rect 73245 587892 73311 587893
rect 73705 587892 73771 587893
rect 71262 587890 71268 587892
rect 69749 587832 69754 587888
rect 68756 587828 68762 587830
rect 69749 587828 69796 587832
rect 69860 587830 69906 587890
rect 71129 587888 71268 587890
rect 71129 587832 71134 587888
rect 71190 587832 71268 587888
rect 71129 587830 71268 587832
rect 69860 587828 69866 587830
rect 68645 587827 68711 587828
rect 69749 587827 69815 587828
rect 71129 587827 71195 587830
rect 71262 587828 71268 587830
rect 71332 587828 71338 587892
rect 72141 587888 72188 587892
rect 72252 587890 72258 587892
rect 72141 587832 72146 587888
rect 72141 587828 72188 587832
rect 72252 587830 72298 587890
rect 73245 587888 73292 587892
rect 73356 587890 73362 587892
rect 73654 587890 73660 587892
rect 73245 587832 73250 587888
rect 72252 587828 72258 587830
rect 73245 587828 73292 587832
rect 73356 587830 73402 587890
rect 73614 587830 73660 587890
rect 73724 587888 73771 587892
rect 73766 587832 73771 587888
rect 73356 587828 73362 587830
rect 73654 587828 73660 587830
rect 73724 587828 73771 587832
rect 72141 587827 72207 587828
rect 73245 587827 73311 587828
rect 73705 587827 73771 587828
rect 74349 587892 74415 587893
rect 76097 587892 76163 587893
rect 74349 587888 74396 587892
rect 74460 587890 74466 587892
rect 76046 587890 76052 587892
rect 74349 587832 74354 587888
rect 74349 587828 74396 587832
rect 74460 587830 74506 587890
rect 76006 587830 76052 587890
rect 76116 587888 76163 587892
rect 76158 587832 76163 587888
rect 74460 587828 74466 587830
rect 76046 587828 76052 587830
rect 76116 587828 76163 587832
rect 74349 587827 74415 587828
rect 76097 587827 76163 587828
rect 77385 587890 77451 587893
rect 78489 587892 78555 587893
rect 78070 587890 78076 587892
rect 77385 587888 78076 587890
rect 77385 587832 77390 587888
rect 77446 587832 78076 587888
rect 77385 587830 78076 587832
rect 77385 587827 77451 587830
rect 78070 587828 78076 587830
rect 78140 587828 78146 587892
rect 78438 587890 78444 587892
rect 78398 587830 78444 587890
rect 78508 587888 78555 587892
rect 78550 587832 78555 587888
rect 78438 587828 78444 587830
rect 78508 587828 78555 587832
rect 78489 587827 78555 587828
rect 79133 587892 79199 587893
rect 81065 587892 81131 587893
rect 83641 587892 83707 587893
rect 88241 587892 88307 587893
rect 91001 587892 91067 587893
rect 93577 587892 93643 587893
rect 79133 587888 79180 587892
rect 79244 587890 79250 587892
rect 81014 587890 81020 587892
rect 79133 587832 79138 587888
rect 79133 587828 79180 587832
rect 79244 587830 79290 587890
rect 80974 587830 81020 587890
rect 81084 587888 81131 587892
rect 83590 587890 83596 587892
rect 81126 587832 81131 587888
rect 79244 587828 79250 587830
rect 81014 587828 81020 587830
rect 81084 587828 81131 587832
rect 83550 587830 83596 587890
rect 83660 587888 83707 587892
rect 88190 587890 88196 587892
rect 83702 587832 83707 587888
rect 83590 587828 83596 587830
rect 83660 587828 83707 587832
rect 88150 587830 88196 587890
rect 88260 587888 88307 587892
rect 90950 587890 90956 587892
rect 88302 587832 88307 587888
rect 88190 587828 88196 587830
rect 88260 587828 88307 587832
rect 90910 587830 90956 587890
rect 91020 587888 91067 587892
rect 93526 587890 93532 587892
rect 91062 587832 91067 587888
rect 90950 587828 90956 587830
rect 91020 587828 91067 587832
rect 93486 587830 93532 587890
rect 93596 587888 93643 587892
rect 93638 587832 93643 587888
rect 93526 587828 93532 587830
rect 93596 587828 93643 587832
rect 95918 587828 95924 587892
rect 95988 587890 95994 587892
rect 96061 587890 96127 587893
rect 98545 587892 98611 587893
rect 100937 587892 101003 587893
rect 98494 587890 98500 587892
rect 95988 587888 96127 587890
rect 95988 587832 96066 587888
rect 96122 587832 96127 587888
rect 95988 587830 96127 587832
rect 98454 587830 98500 587890
rect 98564 587888 98611 587892
rect 100886 587890 100892 587892
rect 98606 587832 98611 587888
rect 95988 587828 95994 587830
rect 79133 587827 79199 587828
rect 81065 587827 81131 587828
rect 83641 587827 83707 587828
rect 88241 587827 88307 587828
rect 91001 587827 91067 587828
rect 93577 587827 93643 587828
rect 96061 587827 96127 587830
rect 98494 587828 98500 587830
rect 98564 587828 98611 587832
rect 100846 587830 100892 587890
rect 100956 587888 101003 587892
rect 100998 587832 101003 587888
rect 100886 587828 100892 587830
rect 100956 587828 101003 587832
rect 103462 587828 103468 587892
rect 103532 587890 103538 587892
rect 103605 587890 103671 587893
rect 103532 587888 103671 587890
rect 103532 587832 103610 587888
rect 103666 587832 103671 587888
rect 103532 587830 103671 587832
rect 103532 587828 103538 587830
rect 98545 587827 98611 587828
rect 100937 587827 101003 587828
rect 103605 587827 103671 587830
rect 105537 587890 105603 587893
rect 108389 587892 108455 587893
rect 105854 587890 105860 587892
rect 105537 587888 105860 587890
rect 105537 587832 105542 587888
rect 105598 587832 105860 587888
rect 105537 587830 105860 587832
rect 105537 587827 105603 587830
rect 105854 587828 105860 587830
rect 105924 587828 105930 587892
rect 108389 587888 108436 587892
rect 108500 587890 108506 587892
rect 108389 587832 108394 587888
rect 108389 587828 108436 587832
rect 108500 587830 108546 587890
rect 108500 587828 108506 587830
rect 111006 587828 111012 587892
rect 111076 587890 111082 587892
rect 111241 587890 111307 587893
rect 111076 587888 111307 587890
rect 111076 587832 111246 587888
rect 111302 587832 111307 587888
rect 111076 587830 111307 587832
rect 111076 587828 111082 587830
rect 108389 587827 108455 587828
rect 111241 587827 111307 587830
rect 113398 587828 113404 587892
rect 113468 587890 113474 587892
rect 113817 587890 113883 587893
rect 113468 587888 113883 587890
rect 113468 587832 113822 587888
rect 113878 587832 113883 587888
rect 113468 587830 113883 587832
rect 113468 587828 113474 587830
rect 113817 587827 113883 587830
rect 114553 587890 114619 587893
rect 115790 587890 115796 587892
rect 114553 587888 115796 587890
rect 114553 587832 114558 587888
rect 114614 587832 115796 587888
rect 114553 587830 115796 587832
rect 114553 587827 114619 587830
rect 115790 587828 115796 587830
rect 115860 587828 115866 587892
rect 118141 587890 118207 587893
rect 118366 587890 118372 587892
rect 118141 587888 118372 587890
rect 118141 587832 118146 587888
rect 118202 587832 118372 587888
rect 118141 587830 118372 587832
rect 118141 587827 118207 587830
rect 118366 587828 118372 587830
rect 118436 587828 118442 587892
rect 120533 587890 120599 587893
rect 125961 587892 126027 587893
rect 120942 587890 120948 587892
rect 120533 587888 120948 587890
rect 120533 587832 120538 587888
rect 120594 587832 120948 587888
rect 120533 587830 120948 587832
rect 120533 587827 120599 587830
rect 120942 587828 120948 587830
rect 121012 587828 121018 587892
rect 125910 587890 125916 587892
rect 125870 587830 125916 587890
rect 125980 587888 126027 587892
rect 126022 587832 126027 587888
rect 125910 587828 125916 587830
rect 125980 587828 126027 587832
rect 125961 587827 126027 587828
rect 436277 587890 436343 587893
rect 438117 587892 438183 587893
rect 439589 587892 439655 587893
rect 441613 587892 441679 587893
rect 443085 587892 443151 587893
rect 444189 587892 444255 587893
rect 437054 587890 437060 587892
rect 436277 587888 437060 587890
rect 436277 587832 436282 587888
rect 436338 587832 437060 587888
rect 436277 587830 437060 587832
rect 436277 587827 436343 587830
rect 437054 587828 437060 587830
rect 437124 587828 437130 587892
rect 438117 587888 438164 587892
rect 438228 587890 438234 587892
rect 438117 587832 438122 587888
rect 438117 587828 438164 587832
rect 438228 587830 438274 587890
rect 439589 587888 439636 587892
rect 439700 587890 439706 587892
rect 439589 587832 439594 587888
rect 438228 587828 438234 587830
rect 439589 587828 439636 587832
rect 439700 587830 439746 587890
rect 441613 587888 441660 587892
rect 441724 587890 441730 587892
rect 441613 587832 441618 587888
rect 439700 587828 439706 587830
rect 441613 587828 441660 587832
rect 441724 587830 441770 587890
rect 443085 587888 443132 587892
rect 443196 587890 443202 587892
rect 443085 587832 443090 587888
rect 441724 587828 441730 587830
rect 443085 587828 443132 587832
rect 443196 587830 443242 587890
rect 444189 587888 444236 587892
rect 444300 587890 444306 587892
rect 444189 587832 444194 587888
rect 443196 587828 443202 587830
rect 444189 587828 444236 587832
rect 444300 587830 444346 587890
rect 444300 587828 444306 587830
rect 445518 587828 445524 587892
rect 445588 587890 445594 587892
rect 445661 587890 445727 587893
rect 446489 587892 446555 587893
rect 446438 587890 446444 587892
rect 445588 587888 445727 587890
rect 445588 587832 445666 587888
rect 445722 587832 445727 587888
rect 445588 587830 445727 587832
rect 446398 587830 446444 587890
rect 446508 587888 446555 587892
rect 446550 587832 446555 587888
rect 445588 587828 445594 587830
rect 438117 587827 438183 587828
rect 439589 587827 439655 587828
rect 441613 587827 441679 587828
rect 443085 587827 443151 587828
rect 444189 587827 444255 587828
rect 445661 587827 445727 587830
rect 446438 587828 446444 587830
rect 446508 587828 446555 587832
rect 446489 587827 446555 587828
rect 447317 587890 447383 587893
rect 447542 587890 447548 587892
rect 447317 587888 447548 587890
rect 447317 587832 447322 587888
rect 447378 587832 447548 587888
rect 447317 587830 447548 587832
rect 447317 587827 447383 587830
rect 447542 587828 447548 587830
rect 447612 587828 447618 587892
rect 448513 587890 448579 587893
rect 449893 587892 449959 587893
rect 450629 587892 450695 587893
rect 453573 587892 453639 587893
rect 454585 587892 454651 587893
rect 448646 587890 448652 587892
rect 448513 587888 448652 587890
rect 448513 587832 448518 587888
rect 448574 587832 448652 587888
rect 448513 587830 448652 587832
rect 448513 587827 448579 587830
rect 448646 587828 448652 587830
rect 448716 587828 448722 587892
rect 449893 587890 449940 587892
rect 449848 587888 449940 587890
rect 449848 587832 449898 587888
rect 449848 587830 449940 587832
rect 449893 587828 449940 587830
rect 450004 587828 450010 587892
rect 450629 587888 450676 587892
rect 450740 587890 450746 587892
rect 450629 587832 450634 587888
rect 450629 587828 450676 587832
rect 450740 587830 450786 587890
rect 453573 587888 453620 587892
rect 453684 587890 453690 587892
rect 454534 587890 454540 587892
rect 453573 587832 453578 587888
rect 450740 587828 450746 587830
rect 453573 587828 453620 587832
rect 453684 587830 453730 587890
rect 454494 587830 454540 587890
rect 454604 587888 454651 587892
rect 454646 587832 454651 587888
rect 453684 587828 453690 587830
rect 454534 587828 454540 587830
rect 454604 587828 454651 587832
rect 449893 587827 449959 587828
rect 450629 587827 450695 587828
rect 453573 587827 453639 587828
rect 454585 587827 454651 587828
rect 456057 587890 456123 587893
rect 456190 587890 456196 587892
rect 456057 587888 456196 587890
rect 456057 587832 456062 587888
rect 456118 587832 456196 587888
rect 456057 587830 456196 587832
rect 456057 587827 456123 587830
rect 456190 587828 456196 587830
rect 456260 587828 456266 587892
rect 456793 587890 456859 587893
rect 456926 587890 456932 587892
rect 456793 587888 456932 587890
rect 456793 587832 456798 587888
rect 456854 587832 456932 587888
rect 456793 587830 456932 587832
rect 456793 587827 456859 587830
rect 456926 587828 456932 587830
rect 456996 587828 457002 587892
rect 457253 587890 457319 587893
rect 471237 587892 471303 587893
rect 472157 587892 472223 587893
rect 473353 587892 473419 587893
rect 458030 587890 458036 587892
rect 457253 587888 458036 587890
rect 457253 587832 457258 587888
rect 457314 587832 458036 587888
rect 457253 587830 458036 587832
rect 457253 587827 457319 587830
rect 458030 587828 458036 587830
rect 458100 587890 458106 587892
rect 458100 587830 470610 587890
rect 458100 587828 458106 587830
rect 19149 587754 19215 587757
rect 48589 587756 48655 587757
rect 50061 587756 50127 587757
rect 35934 587754 35940 587756
rect 19149 587752 35940 587754
rect 19149 587696 19154 587752
rect 19210 587696 35940 587752
rect 19149 587694 35940 587696
rect 19149 587691 19215 587694
rect 35934 587692 35940 587694
rect 36004 587692 36010 587756
rect 48589 587752 48636 587756
rect 48700 587754 48706 587756
rect 48589 587696 48594 587752
rect 48589 587692 48636 587696
rect 48700 587694 48746 587754
rect 50061 587752 50108 587756
rect 50172 587754 50178 587756
rect 52637 587754 52703 587757
rect 53414 587754 53420 587756
rect 50061 587696 50066 587752
rect 48700 587692 48706 587694
rect 50061 587692 50108 587696
rect 50172 587694 50218 587754
rect 52637 587752 53420 587754
rect 52637 587696 52642 587752
rect 52698 587696 53420 587752
rect 52637 587694 53420 587696
rect 50172 587692 50178 587694
rect 48589 587691 48655 587692
rect 50061 587691 50127 587692
rect 52637 587691 52703 587694
rect 53414 587692 53420 587694
rect 53484 587692 53490 587756
rect 59486 587692 59492 587756
rect 59556 587754 59562 587756
rect 59813 587754 59879 587757
rect 59556 587752 59879 587754
rect 59556 587696 59818 587752
rect 59874 587696 59879 587752
rect 59556 587694 59879 587696
rect 59556 587692 59562 587694
rect 59813 587691 59879 587694
rect 65517 587754 65583 587757
rect 452377 587756 452443 587757
rect 453481 587756 453547 587757
rect 65517 587752 74550 587754
rect 65517 587696 65522 587752
rect 65578 587696 74550 587752
rect 65517 587694 74550 587696
rect 65517 587691 65583 587694
rect 19742 587556 19748 587620
rect 19812 587618 19818 587620
rect 38142 587618 38148 587620
rect 19812 587558 38148 587618
rect 19812 587556 19818 587558
rect 38142 587556 38148 587558
rect 38212 587556 38218 587620
rect 58198 587556 58204 587620
rect 58268 587618 58274 587620
rect 74490 587618 74550 587694
rect 418838 587692 418844 587756
rect 418908 587754 418914 587756
rect 448278 587754 448284 587756
rect 418908 587694 448284 587754
rect 418908 587692 418914 587694
rect 448278 587692 448284 587694
rect 448348 587692 448354 587756
rect 452326 587754 452332 587756
rect 452286 587694 452332 587754
rect 452396 587752 452443 587756
rect 453430 587754 453436 587756
rect 452438 587696 452443 587752
rect 452326 587692 452332 587694
rect 452396 587692 452443 587696
rect 453390 587694 453436 587754
rect 453500 587752 453547 587756
rect 453542 587696 453547 587752
rect 453430 587692 453436 587694
rect 453500 587692 453547 587696
rect 455822 587692 455828 587756
rect 455892 587754 455898 587756
rect 456149 587754 456215 587757
rect 455892 587752 456215 587754
rect 455892 587696 456154 587752
rect 456210 587696 456215 587752
rect 455892 587694 456215 587696
rect 455892 587692 455898 587694
rect 452377 587691 452443 587692
rect 453481 587691 453547 587692
rect 456149 587691 456215 587694
rect 458265 587754 458331 587757
rect 460657 587756 460723 587757
rect 459318 587754 459324 587756
rect 458265 587752 459324 587754
rect 458265 587696 458270 587752
rect 458326 587696 459324 587752
rect 458265 587694 459324 587696
rect 458265 587691 458331 587694
rect 459318 587692 459324 587694
rect 459388 587692 459394 587756
rect 460606 587754 460612 587756
rect 460566 587694 460612 587754
rect 460676 587752 460723 587756
rect 460718 587696 460723 587752
rect 460606 587692 460612 587694
rect 460676 587692 460723 587696
rect 460657 587691 460723 587692
rect 460933 587756 460999 587757
rect 460933 587752 460980 587756
rect 461044 587754 461050 587756
rect 461577 587754 461643 587757
rect 461710 587754 461716 587756
rect 460933 587696 460938 587752
rect 460933 587692 460980 587696
rect 461044 587694 461090 587754
rect 461577 587752 461716 587754
rect 461577 587696 461582 587752
rect 461638 587696 461716 587752
rect 461577 587694 461716 587696
rect 461044 587692 461050 587694
rect 460933 587691 460999 587692
rect 461577 587691 461643 587694
rect 461710 587692 461716 587694
rect 461780 587692 461786 587756
rect 462313 587754 462379 587757
rect 463877 587756 463943 587757
rect 463550 587754 463556 587756
rect 462313 587752 463556 587754
rect 462313 587696 462318 587752
rect 462374 587696 463556 587752
rect 462313 587694 463556 587696
rect 462313 587691 462379 587694
rect 463550 587692 463556 587694
rect 463620 587692 463626 587756
rect 463877 587752 463924 587756
rect 463988 587754 463994 587756
rect 465073 587754 465139 587757
rect 466269 587756 466335 587757
rect 467557 587756 467623 587757
rect 468661 587756 468727 587757
rect 469765 587756 469831 587757
rect 465942 587754 465948 587756
rect 463877 587696 463882 587752
rect 463877 587692 463924 587696
rect 463988 587694 464034 587754
rect 465073 587752 465948 587754
rect 465073 587696 465078 587752
rect 465134 587696 465948 587752
rect 465073 587694 465948 587696
rect 463988 587692 463994 587694
rect 463877 587691 463943 587692
rect 465073 587691 465139 587694
rect 465942 587692 465948 587694
rect 466012 587692 466018 587756
rect 466269 587752 466316 587756
rect 466380 587754 466386 587756
rect 466269 587696 466274 587752
rect 466269 587692 466316 587696
rect 466380 587694 466426 587754
rect 467557 587752 467604 587756
rect 467668 587754 467674 587756
rect 467557 587696 467562 587752
rect 466380 587692 466386 587694
rect 467557 587692 467604 587696
rect 467668 587694 467714 587754
rect 468661 587752 468708 587756
rect 468772 587754 468778 587756
rect 468661 587696 468666 587752
rect 467668 587692 467674 587694
rect 468661 587692 468708 587696
rect 468772 587694 468818 587754
rect 469765 587752 469812 587756
rect 469876 587754 469882 587756
rect 470550 587754 470610 587830
rect 471237 587888 471284 587892
rect 471348 587890 471354 587892
rect 471237 587832 471242 587888
rect 471237 587828 471284 587832
rect 471348 587830 471394 587890
rect 472157 587888 472204 587892
rect 472268 587890 472274 587892
rect 473302 587890 473308 587892
rect 472157 587832 472162 587888
rect 471348 587828 471354 587830
rect 472157 587828 472204 587832
rect 472268 587830 472314 587890
rect 473262 587830 473308 587890
rect 473372 587888 473419 587892
rect 473414 587832 473419 587888
rect 472268 587828 472274 587830
rect 473302 587828 473308 587830
rect 473372 587828 473419 587832
rect 471237 587827 471303 587828
rect 472157 587827 472223 587828
rect 473353 587827 473419 587828
rect 473629 587890 473695 587893
rect 476941 587892 477007 587893
rect 478045 587892 478111 587893
rect 479149 587892 479215 587893
rect 474406 587890 474412 587892
rect 473629 587888 474412 587890
rect 473629 587832 473634 587888
rect 473690 587832 474412 587888
rect 473629 587830 474412 587832
rect 473629 587827 473695 587830
rect 474406 587828 474412 587830
rect 474476 587828 474482 587892
rect 476941 587888 476988 587892
rect 477052 587890 477058 587892
rect 476941 587832 476946 587888
rect 476941 587828 476988 587832
rect 477052 587830 477098 587890
rect 478045 587888 478092 587892
rect 478156 587890 478162 587892
rect 478045 587832 478050 587888
rect 477052 587828 477058 587830
rect 478045 587828 478092 587832
rect 478156 587830 478202 587890
rect 479149 587888 479196 587892
rect 479260 587890 479266 587892
rect 480253 587890 480319 587893
rect 480846 587890 480852 587892
rect 479149 587832 479154 587888
rect 478156 587828 478162 587830
rect 479149 587828 479196 587832
rect 479260 587830 479306 587890
rect 480253 587888 480852 587890
rect 480253 587832 480258 587888
rect 480314 587832 480852 587888
rect 480253 587830 480852 587832
rect 479260 587828 479266 587830
rect 476941 587827 477007 587828
rect 478045 587827 478111 587828
rect 479149 587827 479215 587828
rect 480253 587827 480319 587830
rect 480846 587828 480852 587830
rect 480916 587828 480922 587892
rect 483013 587890 483079 587893
rect 483422 587890 483428 587892
rect 483013 587888 483428 587890
rect 483013 587832 483018 587888
rect 483074 587832 483428 587888
rect 483013 587830 483428 587832
rect 483013 587827 483079 587830
rect 483422 587828 483428 587830
rect 483492 587828 483498 587892
rect 485773 587890 485839 587893
rect 485998 587890 486004 587892
rect 485773 587888 486004 587890
rect 485773 587832 485778 587888
rect 485834 587832 486004 587888
rect 485773 587830 486004 587832
rect 485773 587827 485839 587830
rect 485998 587828 486004 587830
rect 486068 587828 486074 587892
rect 487153 587890 487219 587893
rect 488206 587890 488212 587892
rect 487153 587888 488212 587890
rect 487153 587832 487158 587888
rect 487214 587832 488212 587888
rect 487153 587830 488212 587832
rect 487153 587827 487219 587830
rect 488206 587828 488212 587830
rect 488276 587828 488282 587892
rect 492673 587890 492739 587893
rect 493358 587890 493364 587892
rect 492673 587888 493364 587890
rect 492673 587832 492678 587888
rect 492734 587832 493364 587888
rect 492673 587830 493364 587832
rect 492673 587827 492739 587830
rect 493358 587828 493364 587830
rect 493428 587828 493434 587892
rect 495433 587890 495499 587893
rect 495934 587890 495940 587892
rect 495433 587888 495940 587890
rect 495433 587832 495438 587888
rect 495494 587832 495940 587888
rect 495433 587830 495940 587832
rect 495433 587827 495499 587830
rect 495934 587828 495940 587830
rect 496004 587828 496010 587892
rect 498193 587890 498259 587893
rect 500953 587892 501019 587893
rect 498510 587890 498516 587892
rect 498193 587888 498516 587890
rect 498193 587832 498198 587888
rect 498254 587832 498516 587888
rect 498193 587830 498516 587832
rect 498193 587827 498259 587830
rect 498510 587828 498516 587830
rect 498580 587828 498586 587892
rect 500902 587890 500908 587892
rect 500862 587830 500908 587890
rect 500972 587888 501019 587892
rect 501014 587832 501019 587888
rect 500902 587828 500908 587830
rect 500972 587828 501019 587832
rect 500953 587827 501019 587828
rect 502333 587890 502399 587893
rect 503478 587890 503484 587892
rect 502333 587888 503484 587890
rect 502333 587832 502338 587888
rect 502394 587832 503484 587888
rect 502333 587830 503484 587832
rect 502333 587827 502399 587830
rect 503478 587828 503484 587830
rect 503548 587828 503554 587892
rect 505093 587890 505159 587893
rect 505870 587890 505876 587892
rect 505093 587888 505876 587890
rect 505093 587832 505098 587888
rect 505154 587832 505876 587888
rect 505093 587830 505876 587832
rect 505093 587827 505159 587830
rect 505870 587828 505876 587830
rect 505940 587828 505946 587892
rect 507853 587890 507919 587893
rect 508446 587890 508452 587892
rect 507853 587888 508452 587890
rect 507853 587832 507858 587888
rect 507914 587832 508452 587888
rect 507853 587830 508452 587832
rect 507853 587827 507919 587830
rect 508446 587828 508452 587830
rect 508516 587828 508522 587892
rect 510613 587890 510679 587893
rect 513373 587892 513439 587893
rect 511022 587890 511028 587892
rect 510613 587888 511028 587890
rect 510613 587832 510618 587888
rect 510674 587832 511028 587888
rect 510613 587830 511028 587832
rect 510613 587827 510679 587830
rect 511022 587828 511028 587830
rect 511092 587828 511098 587892
rect 513373 587888 513420 587892
rect 513484 587890 513490 587892
rect 514753 587890 514819 587893
rect 515806 587890 515812 587892
rect 513373 587832 513378 587888
rect 513373 587828 513420 587832
rect 513484 587830 513530 587890
rect 514753 587888 515812 587890
rect 514753 587832 514758 587888
rect 514814 587832 515812 587888
rect 514753 587830 515812 587832
rect 513484 587828 513490 587830
rect 513373 587827 513439 587828
rect 514753 587827 514819 587830
rect 515806 587828 515812 587830
rect 515876 587828 515882 587892
rect 517462 587828 517468 587892
rect 517532 587890 517538 587892
rect 518382 587890 518388 587892
rect 517532 587830 518388 587890
rect 517532 587828 517538 587830
rect 518382 587828 518388 587830
rect 518452 587828 518458 587892
rect 520273 587890 520339 587893
rect 523309 587892 523375 587893
rect 525885 587892 525951 587893
rect 520958 587890 520964 587892
rect 520273 587888 520964 587890
rect 520273 587832 520278 587888
rect 520334 587832 520964 587888
rect 520273 587830 520964 587832
rect 520273 587827 520339 587830
rect 520958 587828 520964 587830
rect 521028 587828 521034 587892
rect 523309 587888 523356 587892
rect 523420 587890 523426 587892
rect 523309 587832 523314 587888
rect 523309 587828 523356 587832
rect 523420 587830 523466 587890
rect 525885 587888 525932 587892
rect 525996 587890 526002 587892
rect 525885 587832 525890 587888
rect 523420 587828 523426 587830
rect 525885 587828 525932 587832
rect 525996 587830 526042 587890
rect 525996 587828 526002 587830
rect 523309 587827 523375 587828
rect 525885 587827 525951 587828
rect 473261 587754 473327 587757
rect 469765 587696 469770 587752
rect 468772 587692 468778 587694
rect 469765 587692 469812 587696
rect 469876 587694 469922 587754
rect 470550 587752 473327 587754
rect 470550 587696 473266 587752
rect 473322 587696 473327 587752
rect 470550 587694 473327 587696
rect 469876 587692 469882 587694
rect 466269 587691 466335 587692
rect 467557 587691 467623 587692
rect 468661 587691 468727 587692
rect 469765 587691 469831 587692
rect 473261 587691 473327 587694
rect 75678 587618 75684 587620
rect 58268 587558 70410 587618
rect 74490 587558 75684 587618
rect 58268 587556 58274 587558
rect 57053 587484 57119 587485
rect 19926 587420 19932 587484
rect 19996 587482 20002 587484
rect 40534 587482 40540 587484
rect 19996 587422 40540 587482
rect 19996 587420 20002 587422
rect 40534 587420 40540 587422
rect 40604 587420 40610 587484
rect 57053 587482 57100 587484
rect 56972 587480 57100 587482
rect 57164 587482 57170 587484
rect 65517 587482 65583 587485
rect 65977 587484 66043 587485
rect 65926 587482 65932 587484
rect 57164 587480 65583 587482
rect 56972 587424 57058 587480
rect 57164 587424 65522 587480
rect 65578 587424 65583 587480
rect 56972 587422 57100 587424
rect 57053 587420 57100 587422
rect 57164 587422 65583 587424
rect 65886 587422 65932 587482
rect 65996 587480 66043 587484
rect 66038 587424 66043 587480
rect 57164 587420 57170 587422
rect 57053 587419 57119 587420
rect 65517 587419 65583 587422
rect 65926 587420 65932 587422
rect 65996 587420 66043 587424
rect 68318 587420 68324 587484
rect 68388 587482 68394 587484
rect 68553 587482 68619 587485
rect 68388 587480 68619 587482
rect 68388 587424 68558 587480
rect 68614 587424 68619 587480
rect 68388 587422 68619 587424
rect 70350 587482 70410 587558
rect 75678 587556 75684 587558
rect 75748 587556 75754 587620
rect 419165 587618 419231 587621
rect 473486 587618 473492 587620
rect 419165 587616 473492 587618
rect 419165 587560 419170 587616
rect 419226 587560 473492 587616
rect 419165 587558 473492 587560
rect 419165 587555 419231 587558
rect 473486 587556 473492 587558
rect 473556 587556 473562 587620
rect 76966 587482 76972 587484
rect 70350 587422 76972 587482
rect 68388 587420 68394 587422
rect 65977 587419 66043 587420
rect 68553 587419 68619 587422
rect 76966 587420 76972 587422
rect 77036 587420 77042 587484
rect 418705 587482 418771 587485
rect 476062 587482 476068 587484
rect 418705 587480 476068 587482
rect 418705 587424 418710 587480
rect 418766 587424 476068 587480
rect 418705 587422 476068 587424
rect 418705 587419 418771 587422
rect 476062 587420 476068 587422
rect 476132 587420 476138 587484
rect 19006 587284 19012 587348
rect 19076 587346 19082 587348
rect 41822 587346 41828 587348
rect 19076 587286 41828 587346
rect 19076 587284 19082 587286
rect 41822 587284 41828 587286
rect 41892 587284 41898 587348
rect 61142 587284 61148 587348
rect 61212 587346 61218 587348
rect 61837 587346 61903 587349
rect 61212 587344 61903 587346
rect 61212 587288 61842 587344
rect 61898 587288 61903 587344
rect 61212 587286 61903 587288
rect 61212 587284 61218 587286
rect 61837 587283 61903 587286
rect 63534 587284 63540 587348
rect 63604 587346 63610 587348
rect 63953 587346 64019 587349
rect 63604 587344 64019 587346
rect 63604 587288 63958 587344
rect 64014 587288 64019 587344
rect 63604 587286 64019 587288
rect 63604 587284 63610 587286
rect 63953 587283 64019 587286
rect 85982 587284 85988 587348
rect 86052 587346 86058 587348
rect 195094 587346 195100 587348
rect 86052 587286 195100 587346
rect 86052 587284 86058 587286
rect 195094 587284 195100 587286
rect 195164 587284 195170 587348
rect 418981 587346 419047 587349
rect 478454 587346 478460 587348
rect 418981 587344 478460 587346
rect 418981 587288 418986 587344
rect 419042 587288 478460 587344
rect 418981 587286 478460 587288
rect 418981 587283 419047 587286
rect 478454 587284 478460 587286
rect 478524 587284 478530 587348
rect 16021 587210 16087 587213
rect 58198 587210 58204 587212
rect 16021 587208 58204 587210
rect 16021 587152 16026 587208
rect 16082 587152 58204 587208
rect 16021 587150 58204 587152
rect 16021 587147 16087 587150
rect 58198 587148 58204 587150
rect 58268 587148 58274 587212
rect 70894 587148 70900 587212
rect 70964 587210 70970 587212
rect 198038 587210 198044 587212
rect 70964 587150 198044 587210
rect 70964 587148 70970 587150
rect 198038 587148 198044 587150
rect 198108 587148 198114 587212
rect 388437 587210 388503 587213
rect 458173 587210 458239 587213
rect 462773 587212 462839 587213
rect 465165 587212 465231 587213
rect 458398 587210 458404 587212
rect 388437 587208 451290 587210
rect 388437 587152 388442 587208
rect 388498 587152 451290 587208
rect 388437 587150 451290 587152
rect 388437 587147 388503 587150
rect 122782 587012 122788 587076
rect 122852 587074 122858 587076
rect 122925 587074 122991 587077
rect 122852 587072 122991 587074
rect 122852 587016 122930 587072
rect 122986 587016 122991 587072
rect 122852 587014 122991 587016
rect 122852 587012 122858 587014
rect 122925 587011 122991 587014
rect 419758 587012 419764 587076
rect 419828 587074 419834 587076
rect 436134 587074 436140 587076
rect 419828 587014 436140 587074
rect 419828 587012 419834 587014
rect 436134 587012 436140 587014
rect 436204 587012 436210 587076
rect 451230 587074 451290 587150
rect 458173 587208 458404 587210
rect 458173 587152 458178 587208
rect 458234 587152 458404 587208
rect 458173 587150 458404 587152
rect 458173 587147 458239 587150
rect 458398 587148 458404 587150
rect 458468 587148 458474 587212
rect 462773 587208 462820 587212
rect 462884 587210 462890 587212
rect 462773 587152 462778 587208
rect 462773 587148 462820 587152
rect 462884 587150 462930 587210
rect 465165 587208 465212 587212
rect 465276 587210 465282 587212
rect 465165 587152 465170 587208
rect 462884 587148 462890 587150
rect 465165 587148 465212 587152
rect 465276 587150 465322 587210
rect 465276 587148 465282 587150
rect 462773 587147 462839 587148
rect 465165 587147 465231 587148
rect 468334 587074 468340 587076
rect 451230 587014 468340 587074
rect 468334 587012 468340 587014
rect 468404 587012 468410 587076
rect 417366 586876 417372 586940
rect 417436 586938 417442 586940
rect 417693 586938 417759 586941
rect 417436 586936 417759 586938
rect 417436 586880 417698 586936
rect 417754 586880 417759 586936
rect 417436 586878 417759 586880
rect 417436 586876 417442 586878
rect 417693 586875 417759 586878
rect 451365 586940 451431 586941
rect 451365 586936 451412 586940
rect 451476 586938 451482 586940
rect 456793 586938 456859 586941
rect 475694 586938 475700 586940
rect 451365 586880 451370 586936
rect 451365 586876 451412 586880
rect 451476 586878 451522 586938
rect 456793 586936 475700 586938
rect 456793 586880 456798 586936
rect 456854 586880 475700 586936
rect 456793 586878 475700 586880
rect 451476 586876 451482 586878
rect 451365 586875 451431 586876
rect 456793 586875 456859 586878
rect 475694 586876 475700 586878
rect 475764 586876 475770 586940
rect 417734 586740 417740 586804
rect 417804 586802 417810 586804
rect 440550 586802 440556 586804
rect 417804 586742 440556 586802
rect 417804 586740 417810 586742
rect 440550 586740 440556 586742
rect 440620 586740 440626 586804
rect 470593 586532 470659 586533
rect 489913 586532 489979 586533
rect 470542 586468 470548 586532
rect 470612 586530 470659 586532
rect 470612 586528 470704 586530
rect 470654 586472 470704 586528
rect 470612 586470 470704 586472
rect 470612 586468 470659 586470
rect 489862 586468 489868 586532
rect 489932 586530 489979 586532
rect 489932 586528 490024 586530
rect 489974 586472 490024 586528
rect 489932 586470 490024 586472
rect 489932 586468 489979 586470
rect 470593 586467 470659 586468
rect 489913 586467 489979 586468
rect 157333 585714 157399 585717
rect 199510 585714 199516 585716
rect 157333 585712 199516 585714
rect 157333 585656 157338 585712
rect 157394 585656 199516 585712
rect 157333 585654 199516 585656
rect 157333 585651 157399 585654
rect 199510 585652 199516 585654
rect 199580 585652 199586 585716
rect 376334 585652 376340 585716
rect 376404 585714 376410 585716
rect 517462 585714 517468 585716
rect 376404 585654 517468 585714
rect 376404 585652 376410 585654
rect 517462 585652 517468 585654
rect 517532 585652 517538 585716
rect 150709 585308 150775 585309
rect 550817 585308 550883 585309
rect 150709 585304 150756 585308
rect 150820 585306 150826 585308
rect 550766 585306 550772 585308
rect 150709 585248 150714 585304
rect 150709 585244 150756 585248
rect 150820 585246 150866 585306
rect 550726 585246 550772 585306
rect 550836 585304 550883 585308
rect 550878 585248 550883 585304
rect 150820 585244 150826 585246
rect 550766 585244 550772 585246
rect 550836 585244 550883 585248
rect 150709 585243 150775 585244
rect 550817 585243 550883 585244
rect 419390 584836 419396 584900
rect 419460 584898 419466 584900
rect 436277 584898 436343 584901
rect 419460 584896 436343 584898
rect 419460 584840 436282 584896
rect 436338 584840 436343 584896
rect 419460 584838 436343 584840
rect 419460 584836 419466 584838
rect 436277 584835 436343 584838
rect 378133 584762 378199 584765
rect 379053 584762 379119 584765
rect 378133 584760 379119 584762
rect 378133 584704 378138 584760
rect 378194 584704 379058 584760
rect 379114 584704 379119 584760
rect 378133 584702 379119 584704
rect 378133 584699 378199 584702
rect 379053 584699 379119 584702
rect 413277 584762 413343 584765
rect 460933 584762 460999 584765
rect 413277 584760 460999 584762
rect 413277 584704 413282 584760
rect 413338 584704 460938 584760
rect 460994 584704 460999 584760
rect 413277 584702 460999 584704
rect 413277 584699 413343 584702
rect 460933 584699 460999 584702
rect 122925 584626 122991 584629
rect 197854 584626 197860 584628
rect 122925 584624 197860 584626
rect 122925 584568 122930 584624
rect 122986 584568 197860 584624
rect 122925 584566 197860 584568
rect 122925 584563 122991 584566
rect 197854 584564 197860 584566
rect 197924 584564 197930 584628
rect 379053 584626 379119 584629
rect 465073 584626 465139 584629
rect 379053 584624 465139 584626
rect 379053 584568 379058 584624
rect 379114 584568 465078 584624
rect 465134 584568 465139 584624
rect 379053 584566 465139 584568
rect 379053 584563 379119 584566
rect 465073 584563 465139 584566
rect 120533 584490 120599 584493
rect 201350 584490 201356 584492
rect 120533 584488 201356 584490
rect 120533 584432 120538 584488
rect 120594 584432 201356 584488
rect 120533 584430 201356 584432
rect 120533 584427 120599 584430
rect 201350 584428 201356 584430
rect 201420 584428 201426 584492
rect 377857 584490 377923 584493
rect 507853 584490 507919 584493
rect 377857 584488 507919 584490
rect 377857 584432 377862 584488
rect 377918 584432 507858 584488
rect 507914 584432 507919 584488
rect 377857 584430 507919 584432
rect 377857 584427 377923 584430
rect 507853 584427 507919 584430
rect 118141 584354 118207 584357
rect 199694 584354 199700 584356
rect 118141 584352 199700 584354
rect 118141 584296 118146 584352
rect 118202 584296 199700 584352
rect 118141 584294 199700 584296
rect 118141 584291 118207 584294
rect 199694 584292 199700 584294
rect 199764 584292 199770 584356
rect 374494 584292 374500 584356
rect 374564 584354 374570 584356
rect 514753 584354 514819 584357
rect 374564 584352 514819 584354
rect 374564 584296 514758 584352
rect 514814 584296 514819 584352
rect 374564 584294 514819 584296
rect 374564 584292 374570 584294
rect 514753 584291 514819 584294
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 156558 579186 156618 579190
rect 158713 579186 158779 579189
rect 156558 579184 158779 579186
rect 156558 579128 158718 579184
rect 158774 579128 158779 579184
rect 156558 579126 158779 579128
rect 556570 579186 556630 579190
rect 558913 579186 558979 579189
rect 556570 579184 558979 579186
rect 556570 579128 558918 579184
rect 558974 579128 558979 579184
rect 556570 579126 558979 579128
rect 158713 579123 158779 579126
rect 558913 579123 558979 579126
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 199878 577084 199884 577148
rect 199948 577084 199954 577148
rect 199886 576876 199946 577084
rect 199878 576812 199884 576876
rect 199948 576812 199954 576876
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 19382 536893 20056 536924
rect 17585 536890 17651 536893
rect 19333 536890 20056 536893
rect 17585 536888 20056 536890
rect 17585 536832 17590 536888
rect 17646 536832 19338 536888
rect 19394 536864 20056 536888
rect 417509 536890 417575 536893
rect 419398 536890 420072 536924
rect 417509 536888 420072 536890
rect 19394 536832 19442 536864
rect 17585 536830 19442 536832
rect 417509 536832 417514 536888
rect 417570 536864 420072 536888
rect 417570 536832 419458 536864
rect 417509 536830 419458 536832
rect 17585 536827 17651 536830
rect 19333 536827 19399 536830
rect 417509 536827 417575 536830
rect 17677 535938 17743 535941
rect 19382 535938 20056 535972
rect 17677 535936 20056 535938
rect 17677 535880 17682 535936
rect 17738 535912 20056 535936
rect 417141 535938 417207 535941
rect 419398 535938 420072 535972
rect 417141 535936 420072 535938
rect 17738 535880 19442 535912
rect 17677 535878 19442 535880
rect 417141 535880 417146 535936
rect 417202 535912 420072 535936
rect 417202 535880 419458 535912
rect 417141 535878 419458 535880
rect 17677 535875 17743 535878
rect 417141 535875 417207 535878
rect 16941 533762 17007 533765
rect 17861 533762 17927 533765
rect 19382 533762 20056 533796
rect 16941 533760 20056 533762
rect 16941 533704 16946 533760
rect 17002 533704 17866 533760
rect 17922 533736 20056 533760
rect 417509 533762 417575 533765
rect 418061 533762 418127 533765
rect 419398 533762 420072 533796
rect 417509 533760 420072 533762
rect 17922 533704 19442 533736
rect 16941 533702 19442 533704
rect 417509 533704 417514 533760
rect 417570 533704 418066 533760
rect 418122 533736 420072 533760
rect 418122 533704 419458 533736
rect 417509 533702 419458 533704
rect 16941 533699 17007 533702
rect 17861 533699 17927 533702
rect 417509 533699 417575 533702
rect 418061 533699 418127 533702
rect 407849 533354 407915 533357
rect 407849 533352 412650 533354
rect 407849 533296 407854 533352
rect 407910 533296 412650 533352
rect 407849 533294 412650 533296
rect 407849 533291 407915 533294
rect 412590 532946 412650 533294
rect 417918 532946 417924 532948
rect 412590 532886 417924 532946
rect 417918 532884 417924 532886
rect 417988 532946 417994 532948
rect 417988 532886 419458 532946
rect 417988 532884 417994 532886
rect 419398 532844 419458 532886
rect 17217 532810 17283 532813
rect 17585 532810 17651 532813
rect 19382 532810 20056 532844
rect 17217 532808 20056 532810
rect 17217 532752 17222 532808
rect 17278 532752 17590 532808
rect 17646 532784 20056 532808
rect 419398 532784 420072 532844
rect 17646 532752 19442 532784
rect 17217 532750 19442 532752
rect 17217 532747 17283 532750
rect 17585 532747 17651 532750
rect 17769 531042 17835 531045
rect 19382 531042 20056 531076
rect 17769 531040 20056 531042
rect 17769 530984 17774 531040
rect 17830 531016 20056 531040
rect 416865 531042 416931 531045
rect 417969 531042 418035 531045
rect 419398 531042 420072 531076
rect 416865 531040 420072 531042
rect 17830 530984 19442 531016
rect 17769 530982 19442 530984
rect 416865 530984 416870 531040
rect 416926 530984 417974 531040
rect 418030 531016 420072 531040
rect 418030 530984 419458 531016
rect 416865 530982 419458 530984
rect 17769 530979 17835 530982
rect 416865 530979 416931 530982
rect 417969 530979 418035 530982
rect 18781 529954 18847 529957
rect 19382 529954 20056 529988
rect 18781 529952 20056 529954
rect 18781 529896 18786 529952
rect 18842 529928 20056 529952
rect 416957 529954 417023 529957
rect 419398 529954 420072 529988
rect 416957 529952 420072 529954
rect 18842 529896 19442 529928
rect 18781 529894 19442 529896
rect 416957 529896 416962 529952
rect 417018 529928 420072 529952
rect 417018 529896 419458 529928
rect 416957 529894 419458 529896
rect 18781 529891 18847 529894
rect 416957 529891 417023 529894
rect 17493 528186 17559 528189
rect 19382 528186 20056 528220
rect 17493 528184 20056 528186
rect 17493 528128 17498 528184
rect 17554 528160 20056 528184
rect 17554 528128 19442 528160
rect 17493 528126 19442 528128
rect 17493 528123 17559 528126
rect 417550 528124 417556 528188
rect 417620 528186 417626 528188
rect 419398 528186 420072 528220
rect 417620 528160 420072 528186
rect 417620 528126 419458 528160
rect 417620 528124 417626 528126
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 17493 527234 17559 527237
rect 17902 527234 17908 527236
rect 17493 527232 17908 527234
rect 17493 527176 17498 527232
rect 17554 527176 17908 527232
rect 17493 527174 17908 527176
rect 17493 527171 17559 527174
rect 17902 527172 17908 527174
rect 17972 527172 17978 527236
rect 415853 527234 415919 527237
rect 417550 527234 417556 527236
rect 415853 527232 417556 527234
rect 415853 527176 415858 527232
rect 415914 527176 417556 527232
rect 415853 527174 417556 527176
rect 415853 527171 415919 527174
rect 417550 527172 417556 527174
rect 417620 527172 417626 527236
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 15929 521522 15995 521525
rect 17902 521522 17908 521524
rect 15929 521520 17908 521522
rect 15929 521464 15934 521520
rect 15990 521464 17908 521520
rect 15929 521462 17908 521464
rect 15929 521459 15995 521462
rect 17902 521460 17908 521462
rect 17972 521460 17978 521524
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 19241 509962 19307 509965
rect 19382 509962 20056 509996
rect 19241 509960 20056 509962
rect 19241 509904 19246 509960
rect 19302 509936 20056 509960
rect 416865 509962 416931 509965
rect 417417 509962 417483 509965
rect 419398 509962 420072 509996
rect 416865 509960 420072 509962
rect 19302 509904 19442 509936
rect 19241 509902 19442 509904
rect 416865 509904 416870 509960
rect 416926 509904 417422 509960
rect 417478 509936 420072 509960
rect 417478 509904 419458 509936
rect 416865 509902 419458 509904
rect 19241 509899 19307 509902
rect 416865 509899 416931 509902
rect 417417 509899 417483 509902
rect 16297 508330 16363 508333
rect 19382 508330 20056 508364
rect 16297 508328 20056 508330
rect 16297 508272 16302 508328
rect 16358 508304 20056 508328
rect 417785 508330 417851 508333
rect 419398 508330 420072 508364
rect 417785 508328 420072 508330
rect 16358 508272 19442 508304
rect 16297 508270 19442 508272
rect 417785 508272 417790 508328
rect 417846 508304 420072 508328
rect 417846 508272 419458 508304
rect 417785 508270 419458 508272
rect 16297 508267 16363 508270
rect 417785 508267 417851 508270
rect 19425 508092 19491 508095
rect 19425 508090 20056 508092
rect 19425 508034 19430 508090
rect 19486 508034 20056 508090
rect 19425 508032 20056 508034
rect 417417 508058 417483 508061
rect 419398 508058 420072 508092
rect 417417 508056 420072 508058
rect 19425 508029 19491 508032
rect 417417 508000 417422 508056
rect 417478 508032 420072 508056
rect 417478 508000 419458 508032
rect 417417 507998 419458 508000
rect 417417 507995 417483 507998
rect 199694 505140 199700 505204
rect 199764 505202 199770 505204
rect 200062 505202 200068 505204
rect 199764 505142 200068 505202
rect 199764 505140 199770 505142
rect 200062 505140 200068 505142
rect 200132 505140 200138 505204
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 201125 501666 201191 501669
rect 248454 501666 248460 501668
rect 201125 501664 248460 501666
rect 201125 501608 201130 501664
rect 201186 501608 248460 501664
rect 201125 501606 248460 501608
rect 201125 501603 201191 501606
rect 248454 501604 248460 501606
rect 248524 501604 248530 501668
rect 202454 500788 202460 500852
rect 202524 500850 202530 500852
rect 202524 500790 214114 500850
rect 202524 500788 202530 500790
rect 214054 500717 214114 500790
rect 202270 500652 202276 500716
rect 202340 500714 202346 500716
rect 213913 500714 213979 500717
rect 202340 500712 213979 500714
rect 202340 500656 213918 500712
rect 213974 500656 213979 500712
rect 202340 500654 213979 500656
rect 214054 500712 214163 500717
rect 214054 500656 214102 500712
rect 214158 500656 214163 500712
rect 214054 500654 214163 500656
rect 202340 500652 202346 500654
rect 213913 500651 213979 500654
rect 214097 500651 214163 500654
rect 354857 500714 354923 500717
rect 364149 500714 364215 500717
rect 354857 500712 364215 500714
rect 354857 500656 354862 500712
rect 354918 500656 364154 500712
rect 364210 500656 364215 500712
rect 354857 500654 364215 500656
rect 354857 500651 354923 500654
rect 364149 500651 364215 500654
rect 366357 500714 366423 500717
rect 375414 500714 375420 500716
rect 366357 500712 375420 500714
rect 366357 500656 366362 500712
rect 366418 500656 375420 500712
rect 366357 500654 375420 500656
rect 366357 500651 366423 500654
rect 375414 500652 375420 500654
rect 375484 500652 375490 500716
rect 202086 500516 202092 500580
rect 202156 500578 202162 500580
rect 214005 500578 214071 500581
rect 202156 500576 214071 500578
rect 202156 500520 214010 500576
rect 214066 500520 214071 500576
rect 202156 500518 214071 500520
rect 202156 500516 202162 500518
rect 214005 500515 214071 500518
rect 320173 500578 320239 500581
rect 419165 500578 419231 500581
rect 320173 500576 419231 500578
rect 320173 500520 320178 500576
rect 320234 500520 419170 500576
rect 419226 500520 419231 500576
rect 320173 500518 419231 500520
rect 320173 500515 320239 500518
rect 419165 500515 419231 500518
rect 203374 500380 203380 500444
rect 203444 500442 203450 500444
rect 228449 500442 228515 500445
rect 203444 500440 228515 500442
rect 203444 500384 228454 500440
rect 228510 500384 228515 500440
rect 203444 500382 228515 500384
rect 203444 500380 203450 500382
rect 228449 500379 228515 500382
rect 288433 500442 288499 500445
rect 416037 500442 416103 500445
rect 288433 500440 416103 500442
rect 288433 500384 288438 500440
rect 288494 500384 416042 500440
rect 416098 500384 416103 500440
rect 288433 500382 416103 500384
rect 288433 500379 288499 500382
rect 416037 500379 416103 500382
rect 212533 500306 212599 500309
rect 407757 500306 407823 500309
rect 212533 500304 407823 500306
rect 212533 500248 212538 500304
rect 212594 500248 407762 500304
rect 407818 500248 407823 500304
rect 212533 500246 407823 500248
rect 212533 500243 212599 500246
rect 407757 500243 407823 500246
rect 211153 500170 211219 500173
rect 410517 500170 410583 500173
rect 211153 500168 410583 500170
rect 211153 500112 211158 500168
rect 211214 500112 410522 500168
rect 410578 500112 410583 500168
rect 211153 500110 410583 500112
rect 211153 500107 211219 500110
rect 410517 500107 410583 500110
rect 203190 499972 203196 500036
rect 203260 500034 203266 500036
rect 215293 500034 215359 500037
rect 203260 500032 215359 500034
rect 203260 499976 215298 500032
rect 215354 499976 215359 500032
rect 203260 499974 215359 499976
rect 203260 499972 203266 499974
rect 215293 499971 215359 499974
rect 369117 500034 369183 500037
rect 377765 500034 377831 500037
rect 369117 500032 377831 500034
rect 369117 499976 369122 500032
rect 369178 499976 377770 500032
rect 377826 499976 377831 500032
rect 369117 499974 377831 499976
rect 369117 499971 369183 499974
rect 377765 499971 377831 499974
rect 202638 499836 202644 499900
rect 202708 499898 202714 499900
rect 212625 499898 212691 499901
rect 202708 499896 212691 499898
rect 202708 499840 212630 499896
rect 212686 499840 212691 499896
rect 202708 499838 212691 499840
rect 202708 499836 202714 499838
rect 212625 499835 212691 499838
rect 45369 499628 45435 499629
rect 45369 499624 45438 499628
rect 45369 499568 45374 499624
rect 45430 499568 45438 499624
rect 45369 499564 45438 499568
rect 45502 499626 45508 499628
rect 45502 499566 45526 499626
rect 45502 499564 45508 499566
rect 199694 499564 199700 499628
rect 199764 499626 199770 499628
rect 200062 499626 200068 499628
rect 199764 499566 200068 499626
rect 199764 499564 199770 499566
rect 200062 499564 200068 499566
rect 200132 499564 200138 499628
rect 45369 499563 45435 499564
rect 199510 499428 199516 499492
rect 199580 499490 199586 499492
rect 244917 499490 244983 499493
rect 199580 499488 244983 499490
rect 199580 499432 244922 499488
rect 244978 499432 244983 499488
rect 199580 499430 244983 499432
rect 199580 499428 199586 499430
rect 244917 499427 244983 499430
rect 37273 498130 37339 498133
rect 41873 498132 41939 498133
rect 38142 498130 38148 498132
rect 37273 498128 38148 498130
rect 37273 498072 37278 498128
rect 37334 498072 38148 498128
rect 37273 498070 38148 498072
rect 37273 498067 37339 498070
rect 38142 498068 38148 498070
rect 38212 498068 38218 498132
rect 41822 498130 41828 498132
rect 41782 498070 41828 498130
rect 41892 498128 41939 498132
rect 41934 498072 41939 498128
rect 41822 498068 41828 498070
rect 41892 498068 41939 498072
rect 43110 498068 43116 498132
rect 43180 498130 43186 498132
rect 43437 498130 43503 498133
rect 43180 498128 43503 498130
rect 43180 498072 43442 498128
rect 43498 498072 43503 498128
rect 43180 498070 43503 498072
rect 43180 498068 43186 498070
rect 41873 498067 41939 498068
rect 43437 498067 43503 498070
rect 46606 498068 46612 498132
rect 46676 498130 46682 498132
rect 46841 498130 46907 498133
rect 47577 498132 47643 498133
rect 48681 498132 48747 498133
rect 51441 498132 51507 498133
rect 47526 498130 47532 498132
rect 46676 498128 46907 498130
rect 46676 498072 46846 498128
rect 46902 498072 46907 498128
rect 46676 498070 46907 498072
rect 47486 498070 47532 498130
rect 47596 498128 47643 498132
rect 48630 498130 48636 498132
rect 47638 498072 47643 498128
rect 46676 498068 46682 498070
rect 46841 498067 46907 498070
rect 47526 498068 47532 498070
rect 47596 498068 47643 498072
rect 48590 498070 48636 498130
rect 48700 498128 48747 498132
rect 51390 498130 51396 498132
rect 48742 498072 48747 498128
rect 48630 498068 48636 498070
rect 48700 498068 48747 498072
rect 51350 498070 51396 498130
rect 51460 498128 51507 498132
rect 51502 498072 51507 498128
rect 51390 498068 51396 498070
rect 51460 498068 51507 498072
rect 47577 498067 47643 498068
rect 48681 498067 48747 498068
rect 51441 498067 51507 498068
rect 52177 498130 52243 498133
rect 53465 498132 53531 498133
rect 52310 498130 52316 498132
rect 52177 498128 52316 498130
rect 52177 498072 52182 498128
rect 52238 498072 52316 498128
rect 52177 498070 52316 498072
rect 52177 498067 52243 498070
rect 52310 498068 52316 498070
rect 52380 498068 52386 498132
rect 53414 498130 53420 498132
rect 53374 498070 53420 498130
rect 53484 498128 53531 498132
rect 53526 498072 53531 498128
rect 53414 498068 53420 498070
rect 53484 498068 53531 498072
rect 53465 498067 53531 498068
rect 53833 498130 53899 498133
rect 55857 498132 55923 498133
rect 59537 498132 59603 498133
rect 60641 498132 60707 498133
rect 54518 498130 54524 498132
rect 53833 498128 54524 498130
rect 53833 498072 53838 498128
rect 53894 498072 54524 498128
rect 53833 498070 54524 498072
rect 53833 498067 53899 498070
rect 54518 498068 54524 498070
rect 54588 498068 54594 498132
rect 55806 498130 55812 498132
rect 55766 498070 55812 498130
rect 55876 498128 55923 498132
rect 59486 498130 59492 498132
rect 55918 498072 55923 498128
rect 55806 498068 55812 498070
rect 55876 498068 55923 498072
rect 59446 498070 59492 498130
rect 59556 498128 59603 498132
rect 60590 498130 60596 498132
rect 59598 498072 59603 498128
rect 59486 498068 59492 498070
rect 59556 498068 59603 498072
rect 60550 498070 60596 498130
rect 60660 498128 60707 498132
rect 60702 498072 60707 498128
rect 60590 498068 60596 498070
rect 60660 498068 60707 498072
rect 63534 498068 63540 498132
rect 63604 498130 63610 498132
rect 63677 498130 63743 498133
rect 63604 498128 63743 498130
rect 63604 498072 63682 498128
rect 63738 498072 63743 498128
rect 63604 498070 63743 498072
rect 63604 498068 63610 498070
rect 55857 498067 55923 498068
rect 59537 498067 59603 498068
rect 60641 498067 60707 498068
rect 63677 498067 63743 498070
rect 63902 498068 63908 498132
rect 63972 498130 63978 498132
rect 64137 498130 64203 498133
rect 67633 498132 67699 498133
rect 67582 498130 67588 498132
rect 63972 498128 64203 498130
rect 63972 498072 64142 498128
rect 64198 498072 64203 498128
rect 63972 498070 64203 498072
rect 67542 498070 67588 498130
rect 67652 498128 67699 498132
rect 67694 498072 67699 498128
rect 63972 498068 63978 498070
rect 64137 498067 64203 498070
rect 67582 498068 67588 498070
rect 67652 498068 67699 498072
rect 67633 498067 67699 498068
rect 71221 498132 71287 498133
rect 71221 498128 71268 498132
rect 71332 498130 71338 498132
rect 71957 498130 72023 498133
rect 73705 498132 73771 498133
rect 72182 498130 72188 498132
rect 71221 498072 71226 498128
rect 71221 498068 71268 498072
rect 71332 498070 71378 498130
rect 71957 498128 72188 498130
rect 71957 498072 71962 498128
rect 72018 498072 72188 498128
rect 71957 498070 72188 498072
rect 71332 498068 71338 498070
rect 71221 498067 71287 498068
rect 71957 498067 72023 498070
rect 72182 498068 72188 498070
rect 72252 498068 72258 498132
rect 73654 498130 73660 498132
rect 73614 498070 73660 498130
rect 73724 498128 73771 498132
rect 73766 498072 73771 498128
rect 73654 498068 73660 498070
rect 73724 498068 73771 498072
rect 73705 498067 73771 498068
rect 73981 498130 74047 498133
rect 78121 498132 78187 498133
rect 74390 498130 74396 498132
rect 73981 498128 74396 498130
rect 73981 498072 73986 498128
rect 74042 498072 74396 498128
rect 73981 498070 74396 498072
rect 73981 498067 74047 498070
rect 74390 498068 74396 498070
rect 74460 498068 74466 498132
rect 78070 498130 78076 498132
rect 78030 498070 78076 498130
rect 78140 498128 78187 498132
rect 78182 498072 78187 498128
rect 78070 498068 78076 498070
rect 78140 498068 78187 498072
rect 113398 498068 113404 498132
rect 113468 498130 113474 498132
rect 114461 498130 114527 498133
rect 113468 498128 114527 498130
rect 113468 498072 114466 498128
rect 114522 498072 114527 498128
rect 113468 498070 114527 498072
rect 113468 498068 113474 498070
rect 78121 498067 78187 498068
rect 114461 498067 114527 498070
rect 120942 498068 120948 498132
rect 121012 498130 121018 498132
rect 121361 498130 121427 498133
rect 121012 498128 121427 498130
rect 121012 498072 121366 498128
rect 121422 498072 121427 498128
rect 121012 498070 121427 498072
rect 121012 498068 121018 498070
rect 121361 498067 121427 498070
rect 195421 498130 195487 498133
rect 237649 498130 237715 498133
rect 441613 498132 441679 498133
rect 445293 498132 445359 498133
rect 195421 498128 237715 498130
rect 195421 498072 195426 498128
rect 195482 498072 237654 498128
rect 237710 498072 237715 498128
rect 195421 498070 237715 498072
rect 195421 498067 195487 498070
rect 237649 498067 237715 498070
rect 417734 498068 417740 498132
rect 417804 498130 417810 498132
rect 440550 498130 440556 498132
rect 417804 498070 440556 498130
rect 417804 498068 417810 498070
rect 440550 498068 440556 498070
rect 440620 498068 440626 498132
rect 441613 498128 441660 498132
rect 441724 498130 441730 498132
rect 441613 498072 441618 498128
rect 441613 498068 441660 498072
rect 441724 498070 441770 498130
rect 445293 498128 445340 498132
rect 445404 498130 445410 498132
rect 445293 498072 445298 498128
rect 441724 498068 441730 498070
rect 445293 498068 445340 498072
rect 445404 498070 445450 498130
rect 445404 498068 445410 498070
rect 448646 498068 448652 498132
rect 448716 498130 448722 498132
rect 449157 498130 449223 498133
rect 448716 498128 449223 498130
rect 448716 498072 449162 498128
rect 449218 498072 449223 498128
rect 448716 498070 449223 498072
rect 448716 498068 448722 498070
rect 441613 498067 441679 498068
rect 445293 498067 445359 498068
rect 449157 498067 449223 498070
rect 451038 498068 451044 498132
rect 451108 498130 451114 498132
rect 451273 498130 451339 498133
rect 452377 498132 452443 498133
rect 454585 498132 454651 498133
rect 452326 498130 452332 498132
rect 451108 498128 451339 498130
rect 451108 498072 451278 498128
rect 451334 498072 451339 498128
rect 451108 498070 451339 498072
rect 452286 498070 452332 498130
rect 452396 498128 452443 498132
rect 454534 498130 454540 498132
rect 452438 498072 452443 498128
rect 451108 498068 451114 498070
rect 451273 498067 451339 498070
rect 452326 498068 452332 498070
rect 452396 498068 452443 498072
rect 454494 498070 454540 498130
rect 454604 498128 454651 498132
rect 454646 498072 454651 498128
rect 454534 498068 454540 498070
rect 454604 498068 454651 498072
rect 452377 498067 452443 498068
rect 454585 498067 454651 498068
rect 455505 498130 455571 498133
rect 456190 498130 456196 498132
rect 455505 498128 456196 498130
rect 455505 498072 455510 498128
rect 455566 498072 456196 498128
rect 455505 498070 456196 498072
rect 455505 498067 455571 498070
rect 456190 498068 456196 498070
rect 456260 498068 456266 498132
rect 469213 498130 469279 498133
rect 473353 498132 473419 498133
rect 469806 498130 469812 498132
rect 469213 498128 469812 498130
rect 469213 498072 469218 498128
rect 469274 498072 469812 498128
rect 469213 498070 469812 498072
rect 469213 498067 469279 498070
rect 469806 498068 469812 498070
rect 469876 498068 469882 498132
rect 473302 498068 473308 498132
rect 473372 498130 473419 498132
rect 473537 498130 473603 498133
rect 473670 498130 473676 498132
rect 473372 498128 473464 498130
rect 473414 498072 473464 498128
rect 473372 498070 473464 498072
rect 473537 498128 473676 498130
rect 473537 498072 473542 498128
rect 473598 498072 473676 498128
rect 473537 498070 473676 498072
rect 473372 498068 473419 498070
rect 473353 498067 473419 498068
rect 473537 498067 473603 498070
rect 473670 498068 473676 498070
rect 473740 498068 473746 498132
rect 480529 498130 480595 498133
rect 480846 498130 480852 498132
rect 480529 498128 480852 498130
rect 480529 498072 480534 498128
rect 480590 498072 480852 498128
rect 480529 498070 480852 498072
rect 480529 498067 480595 498070
rect 480846 498068 480852 498070
rect 480916 498068 480922 498132
rect 494697 498130 494763 498133
rect 495934 498130 495940 498132
rect 494697 498128 495940 498130
rect 494697 498072 494702 498128
rect 494758 498072 495940 498128
rect 494697 498070 495940 498072
rect 494697 498067 494763 498070
rect 495934 498068 495940 498070
rect 496004 498068 496010 498132
rect 504357 498130 504423 498133
rect 505870 498130 505876 498132
rect 504357 498128 505876 498130
rect 504357 498072 504362 498128
rect 504418 498072 505876 498128
rect 504357 498070 505876 498072
rect 504357 498067 504423 498070
rect 505870 498068 505876 498070
rect 505940 498068 505946 498132
rect 512637 498130 512703 498133
rect 513414 498130 513420 498132
rect 512637 498128 513420 498130
rect 512637 498072 512642 498128
rect 512698 498072 513420 498128
rect 512637 498070 513420 498072
rect 512637 498067 512703 498070
rect 513414 498068 513420 498070
rect 513484 498068 513490 498132
rect 519537 498130 519603 498133
rect 520958 498130 520964 498132
rect 519537 498128 520964 498130
rect 519537 498072 519542 498128
rect 519598 498072 520964 498128
rect 519537 498070 520964 498072
rect 519537 498067 519603 498070
rect 520958 498068 520964 498070
rect 521028 498068 521034 498132
rect 44173 497996 44239 497997
rect 58157 497996 58223 497997
rect 44173 497992 44220 497996
rect 44284 497994 44290 497996
rect 58157 497994 58204 497996
rect 44173 497936 44178 497992
rect 44173 497932 44220 497936
rect 44284 497934 44330 497994
rect 58076 497992 58204 497994
rect 58268 497994 58274 497996
rect 76557 497994 76623 497997
rect 76966 497994 76972 497996
rect 58268 497992 76972 497994
rect 58076 497936 58162 497992
rect 58268 497936 76562 497992
rect 76618 497936 76972 497992
rect 58076 497934 58204 497936
rect 44284 497932 44290 497934
rect 58157 497932 58204 497934
rect 58268 497934 76972 497936
rect 58268 497932 58274 497934
rect 44173 497931 44239 497932
rect 58157 497931 58223 497932
rect 76557 497931 76623 497934
rect 76966 497932 76972 497934
rect 77036 497932 77042 497996
rect 195830 497932 195836 497996
rect 195900 497994 195906 497996
rect 238937 497994 239003 497997
rect 195900 497992 239003 497994
rect 195900 497936 238942 497992
rect 238998 497936 239003 497992
rect 195900 497934 239003 497936
rect 195900 497932 195906 497934
rect 238937 497931 239003 497934
rect 419390 497932 419396 497996
rect 419460 497994 419466 497996
rect 436185 497994 436251 497997
rect 419460 497992 436251 497994
rect 419460 497936 436190 497992
rect 436246 497936 436251 497992
rect 419460 497934 436251 497936
rect 419460 497932 419466 497934
rect 436185 497931 436251 497934
rect 463693 497994 463759 497997
rect 463918 497994 463924 497996
rect 463693 497992 463924 497994
rect 463693 497936 463698 497992
rect 463754 497936 463924 497992
rect 463693 497934 463924 497936
rect 463693 497931 463759 497934
rect 463918 497932 463924 497934
rect 463988 497932 463994 497996
rect 467833 497994 467899 497997
rect 468702 497994 468708 497996
rect 467833 497992 468708 497994
rect 467833 497936 467838 497992
rect 467894 497936 468708 497992
rect 467833 497934 468708 497936
rect 467833 497931 467899 497934
rect 468702 497932 468708 497934
rect 468772 497932 468778 497996
rect 36169 497860 36235 497861
rect 36118 497858 36124 497860
rect 36078 497798 36124 497858
rect 36188 497856 36235 497860
rect 36230 497800 36235 497856
rect 36118 497796 36124 497798
rect 36188 497796 36235 497800
rect 36169 497795 36235 497796
rect 37181 497860 37247 497861
rect 37181 497856 37228 497860
rect 37292 497858 37298 497860
rect 37181 497800 37186 497856
rect 37181 497796 37228 497800
rect 37292 497798 37338 497858
rect 37292 497796 37298 497798
rect 50102 497796 50108 497860
rect 50172 497858 50178 497860
rect 50245 497858 50311 497861
rect 57053 497860 57119 497861
rect 57053 497858 57100 497860
rect 50172 497856 50311 497858
rect 50172 497800 50250 497856
rect 50306 497800 50311 497856
rect 50172 497798 50311 497800
rect 56972 497856 57100 497858
rect 57164 497858 57170 497860
rect 75177 497858 75243 497861
rect 75678 497858 75684 497860
rect 57164 497856 75684 497858
rect 56972 497800 57058 497856
rect 57164 497800 75182 497856
rect 75238 497800 75684 497856
rect 56972 497798 57100 497800
rect 50172 497796 50178 497798
rect 37181 497795 37247 497796
rect 50245 497795 50311 497798
rect 57053 497796 57100 497798
rect 57164 497798 75684 497800
rect 57164 497796 57170 497798
rect 57053 497795 57119 497796
rect 75177 497795 75243 497798
rect 75678 497796 75684 497798
rect 75748 497796 75754 497860
rect 199878 497796 199884 497860
rect 199948 497858 199954 497860
rect 247033 497858 247099 497861
rect 199948 497856 247099 497858
rect 199948 497800 247038 497856
rect 247094 497800 247099 497856
rect 199948 497798 247099 497800
rect 199948 497796 199954 497798
rect 247033 497795 247099 497798
rect 460565 497860 460631 497861
rect 460565 497856 460612 497860
rect 460676 497858 460682 497860
rect 462313 497858 462379 497861
rect 462814 497858 462820 497860
rect 460565 497800 460570 497856
rect 460565 497796 460612 497800
rect 460676 497798 460722 497858
rect 462313 497856 462820 497858
rect 462313 497800 462318 497856
rect 462374 497800 462820 497856
rect 462313 497798 462820 497800
rect 460676 497796 460682 497798
rect 460565 497795 460631 497796
rect 462313 497795 462379 497798
rect 462814 497796 462820 497798
rect 462884 497796 462890 497860
rect 583520 497844 584960 498084
rect 73153 497722 73219 497725
rect 73286 497722 73292 497724
rect 73153 497720 73292 497722
rect 73153 497664 73158 497720
rect 73214 497664 73292 497720
rect 73153 497662 73292 497664
rect 73153 497659 73219 497662
rect 73286 497660 73292 497662
rect 73356 497660 73362 497724
rect 198457 497722 198523 497725
rect 245653 497722 245719 497725
rect 198457 497720 245719 497722
rect 198457 497664 198462 497720
rect 198518 497664 245658 497720
rect 245714 497664 245719 497720
rect 198457 497662 245719 497664
rect 198457 497659 198523 497662
rect 245653 497659 245719 497662
rect 470869 497722 470935 497725
rect 471278 497722 471284 497724
rect 470869 497720 471284 497722
rect 470869 497664 470874 497720
rect 470930 497664 471284 497720
rect 470869 497662 471284 497664
rect 470869 497659 470935 497662
rect 471278 497660 471284 497662
rect 471348 497660 471354 497724
rect 474733 497722 474799 497725
rect 475694 497722 475700 497724
rect 474733 497720 475700 497722
rect 474733 497664 474738 497720
rect 474794 497664 475700 497720
rect 474733 497662 475700 497664
rect 474733 497659 474799 497662
rect 475694 497660 475700 497662
rect 475764 497660 475770 497724
rect 476113 497722 476179 497725
rect 476982 497722 476988 497724
rect 476113 497720 476988 497722
rect 476113 497664 476118 497720
rect 476174 497664 476988 497720
rect 476113 497662 476988 497664
rect 476113 497659 476179 497662
rect 476982 497660 476988 497662
rect 477052 497660 477058 497724
rect 19926 497524 19932 497588
rect 19996 497586 20002 497588
rect 22093 497586 22159 497589
rect 19996 497584 22159 497586
rect 19996 497528 22098 497584
rect 22154 497528 22159 497584
rect 19996 497526 22159 497528
rect 19996 497524 20002 497526
rect 22093 497523 22159 497526
rect 234705 497586 234771 497589
rect 378174 497586 378180 497588
rect 234705 497584 378180 497586
rect 234705 497528 234710 497584
rect 234766 497528 378180 497584
rect 234705 497526 378180 497528
rect 234705 497523 234771 497526
rect 378174 497524 378180 497526
rect 378244 497524 378250 497588
rect 211245 497450 211311 497453
rect 391197 497450 391263 497453
rect 211245 497448 391263 497450
rect 211245 497392 211250 497448
rect 211306 497392 391202 497448
rect 391258 497392 391263 497448
rect 211245 497390 391263 497392
rect 211245 497387 211311 497390
rect 391197 497387 391263 497390
rect 444189 497452 444255 497453
rect 444189 497448 444236 497452
rect 444300 497450 444306 497452
rect 444189 497392 444194 497448
rect 444189 497388 444236 497392
rect 444300 497390 444346 497450
rect 444300 497388 444306 497390
rect 450118 497388 450124 497452
rect 450188 497450 450194 497452
rect 450537 497450 450603 497453
rect 450188 497448 450603 497450
rect 450188 497392 450542 497448
rect 450598 497392 450603 497448
rect 450188 497390 450603 497392
rect 450188 497388 450194 497390
rect 444189 497387 444255 497388
rect 450537 497387 450603 497390
rect 457437 497450 457503 497453
rect 458030 497450 458036 497452
rect 457437 497448 458036 497450
rect 457437 497392 457442 497448
rect 457498 497392 458036 497448
rect 457437 497390 458036 497392
rect 457437 497387 457503 497390
rect 458030 497388 458036 497390
rect 458100 497450 458106 497452
rect 462497 497450 462563 497453
rect 458100 497448 462563 497450
rect 458100 497392 462502 497448
rect 462558 497392 462563 497448
rect 458100 497390 462563 497392
rect 458100 497388 458106 497390
rect 462497 497387 462563 497390
rect 466453 497450 466519 497453
rect 467598 497450 467604 497452
rect 466453 497448 467604 497450
rect 466453 497392 466458 497448
rect 466514 497392 467604 497448
rect 466453 497390 467604 497392
rect 466453 497387 466519 497390
rect 467598 497388 467604 497390
rect 467668 497388 467674 497452
rect 461117 497314 461183 497317
rect 461710 497314 461716 497316
rect 461117 497312 461716 497314
rect 461117 497256 461122 497312
rect 461178 497256 461716 497312
rect 461117 497254 461716 497256
rect 461117 497251 461183 497254
rect 461710 497252 461716 497254
rect 461780 497252 461786 497316
rect 465073 497314 465139 497317
rect 466310 497314 466316 497316
rect 465073 497312 466316 497314
rect 465073 497256 465078 497312
rect 465134 497256 466316 497312
rect 465073 497254 466316 497256
rect 465073 497251 465139 497254
rect 466310 497252 466316 497254
rect 466380 497252 466386 497316
rect 478873 497314 478939 497317
rect 479190 497314 479196 497316
rect 478873 497312 479196 497314
rect 478873 497256 478878 497312
rect 478934 497256 479196 497312
rect 478873 497254 479196 497256
rect 478873 497251 478939 497254
rect 479190 497252 479196 497254
rect 479260 497252 479266 497316
rect 68277 497178 68343 497181
rect 106089 497180 106155 497181
rect 446673 497180 446739 497181
rect 68686 497178 68692 497180
rect 68277 497176 68692 497178
rect 68277 497120 68282 497176
rect 68338 497120 68692 497176
rect 68277 497118 68692 497120
rect 68277 497115 68343 497118
rect 68686 497116 68692 497118
rect 68756 497116 68762 497180
rect 106038 497178 106044 497180
rect 105998 497118 106044 497178
rect 106108 497176 106155 497180
rect 446622 497178 446628 497180
rect 106150 497120 106155 497176
rect 106038 497116 106044 497118
rect 106108 497116 106155 497120
rect 446582 497118 446628 497178
rect 446692 497176 446739 497180
rect 446734 497120 446739 497176
rect 446622 497116 446628 497118
rect 446692 497116 446739 497120
rect 106089 497115 106155 497116
rect 446673 497115 446739 497116
rect 465073 497178 465139 497181
rect 465206 497178 465212 497180
rect 465073 497176 465212 497178
rect 465073 497120 465078 497176
rect 465134 497120 465212 497176
rect 465073 497118 465212 497120
rect 465073 497115 465139 497118
rect 465206 497116 465212 497118
rect 465276 497116 465282 497180
rect 473353 497178 473419 497181
rect 474406 497178 474412 497180
rect 473353 497176 474412 497178
rect 473353 497120 473358 497176
rect 473414 497120 474412 497176
rect 473353 497118 474412 497120
rect 473353 497115 473419 497118
rect 474406 497116 474412 497118
rect 474476 497116 474482 497180
rect 39665 497044 39731 497045
rect 39614 497042 39620 497044
rect 39574 496982 39620 497042
rect 39684 497040 39731 497044
rect 39726 496984 39731 497040
rect 39614 496980 39620 496982
rect 39684 496980 39731 496984
rect 61694 496980 61700 497044
rect 61764 497042 61770 497044
rect 61837 497042 61903 497045
rect 61764 497040 61903 497042
rect 61764 496984 61842 497040
rect 61898 496984 61903 497040
rect 61764 496982 61903 496984
rect 61764 496980 61770 496982
rect 39665 496979 39731 496980
rect 61837 496979 61903 496982
rect 66253 497044 66319 497045
rect 66253 497040 66300 497044
rect 66364 497042 66370 497044
rect 436185 497042 436251 497045
rect 447777 497044 447843 497045
rect 437054 497042 437060 497044
rect 66253 496984 66258 497040
rect 66253 496980 66300 496984
rect 66364 496982 66410 497042
rect 436185 497040 437060 497042
rect 436185 496984 436190 497040
rect 436246 496984 437060 497040
rect 436185 496982 437060 496984
rect 66364 496980 66370 496982
rect 66253 496979 66319 496980
rect 436185 496979 436251 496982
rect 437054 496980 437060 496982
rect 437124 496980 437130 497044
rect 447726 497042 447732 497044
rect 447686 496982 447732 497042
rect 447796 497040 447843 497044
rect 447838 496984 447843 497040
rect 447726 496980 447732 496982
rect 447796 496980 447843 496984
rect 447777 496979 447843 496980
rect 453297 497042 453363 497045
rect 453430 497042 453436 497044
rect 453297 497040 453436 497042
rect 453297 496984 453302 497040
rect 453358 496984 453436 497040
rect 453297 496982 453436 496984
rect 453297 496979 453363 496982
rect 453430 496980 453436 496982
rect 453500 496980 453506 497044
rect 462037 497042 462103 497045
rect 456934 497040 462103 497042
rect 456934 496984 462042 497040
rect 462098 496984 462103 497040
rect 456934 496982 462103 496984
rect 456934 496909 456994 496982
rect 462037 496979 462103 496982
rect 471973 497042 472039 497045
rect 472198 497042 472204 497044
rect 471973 497040 472204 497042
rect 471973 496984 471978 497040
rect 472034 496984 472204 497040
rect 471973 496982 472204 496984
rect 471973 496979 472039 496982
rect 472198 496980 472204 496982
rect 472268 496980 472274 497044
rect 477585 497042 477651 497045
rect 478454 497042 478460 497044
rect 477585 497040 478460 497042
rect 477585 496984 477590 497040
rect 477646 496984 478460 497040
rect 477585 496982 478460 496984
rect 477585 496979 477651 496982
rect 478454 496980 478460 496982
rect 478524 496980 478530 497044
rect 40585 496908 40651 496909
rect 48313 496908 48379 496909
rect 40534 496906 40540 496908
rect 40494 496846 40540 496906
rect 40604 496904 40651 496908
rect 48262 496906 48268 496908
rect 40646 496848 40651 496904
rect 40534 496844 40540 496846
rect 40604 496844 40651 496848
rect 48222 496846 48268 496906
rect 48332 496904 48379 496908
rect 48374 496848 48379 496904
rect 48262 496844 48268 496846
rect 48332 496844 48379 496848
rect 50838 496844 50844 496908
rect 50908 496906 50914 496908
rect 50981 496906 51047 496909
rect 50908 496904 51047 496906
rect 50908 496848 50986 496904
rect 51042 496848 51047 496904
rect 50908 496846 51047 496848
rect 50908 496844 50914 496846
rect 40585 496843 40651 496844
rect 48313 496843 48379 496844
rect 50981 496843 51047 496846
rect 53598 496844 53604 496908
rect 53668 496906 53674 496908
rect 53741 496906 53807 496909
rect 53668 496904 53807 496906
rect 53668 496848 53746 496904
rect 53802 496848 53807 496904
rect 53668 496846 53807 496848
rect 53668 496844 53674 496846
rect 53741 496843 53807 496846
rect 56174 496844 56180 496908
rect 56244 496906 56250 496908
rect 56501 496906 56567 496909
rect 56244 496904 56567 496906
rect 56244 496848 56506 496904
rect 56562 496848 56567 496904
rect 56244 496846 56567 496848
rect 56244 496844 56250 496846
rect 56501 496843 56567 496846
rect 58566 496844 58572 496908
rect 58636 496906 58642 496908
rect 59261 496906 59327 496909
rect 58636 496904 59327 496906
rect 58636 496848 59266 496904
rect 59322 496848 59327 496904
rect 58636 496846 59327 496848
rect 58636 496844 58642 496846
rect 59261 496843 59327 496846
rect 61142 496844 61148 496908
rect 61212 496906 61218 496908
rect 62021 496906 62087 496909
rect 61212 496904 62087 496906
rect 61212 496848 62026 496904
rect 62082 496848 62087 496904
rect 61212 496846 62087 496848
rect 61212 496844 61218 496846
rect 62021 496843 62087 496846
rect 62757 496908 62823 496909
rect 62757 496904 62804 496908
rect 62868 496906 62874 496908
rect 62757 496848 62762 496904
rect 62757 496844 62804 496848
rect 62868 496846 62914 496906
rect 62868 496844 62874 496846
rect 65374 496844 65380 496908
rect 65444 496906 65450 496908
rect 65517 496906 65583 496909
rect 65444 496904 65583 496906
rect 65444 496848 65522 496904
rect 65578 496848 65583 496904
rect 65444 496846 65583 496848
rect 65444 496844 65450 496846
rect 62757 496843 62823 496844
rect 65517 496843 65583 496846
rect 65926 496844 65932 496908
rect 65996 496906 66002 496908
rect 66161 496906 66227 496909
rect 65996 496904 66227 496906
rect 65996 496848 66166 496904
rect 66222 496848 66227 496904
rect 65996 496846 66227 496848
rect 65996 496844 66002 496846
rect 66161 496843 66227 496846
rect 68318 496844 68324 496908
rect 68388 496906 68394 496908
rect 68553 496906 68619 496909
rect 68388 496904 68619 496906
rect 68388 496848 68558 496904
rect 68614 496848 68619 496904
rect 68388 496846 68619 496848
rect 68388 496844 68394 496846
rect 68553 496843 68619 496846
rect 69657 496906 69723 496909
rect 69790 496906 69796 496908
rect 69657 496904 69796 496906
rect 69657 496848 69662 496904
rect 69718 496848 69796 496904
rect 69657 496846 69796 496848
rect 69657 496843 69723 496846
rect 69790 496844 69796 496846
rect 69860 496844 69866 496908
rect 70894 496844 70900 496908
rect 70964 496906 70970 496908
rect 71681 496906 71747 496909
rect 70964 496904 71747 496906
rect 70964 496848 71686 496904
rect 71742 496848 71747 496904
rect 70964 496846 71747 496848
rect 70964 496844 70970 496846
rect 71681 496843 71747 496846
rect 73286 496844 73292 496908
rect 73356 496906 73362 496908
rect 73797 496906 73863 496909
rect 73356 496904 73863 496906
rect 73356 496848 73802 496904
rect 73858 496848 73863 496904
rect 73356 496846 73863 496848
rect 73356 496844 73362 496846
rect 73797 496843 73863 496846
rect 76046 496844 76052 496908
rect 76116 496906 76122 496908
rect 76833 496906 76899 496909
rect 76116 496904 76899 496906
rect 76116 496848 76838 496904
rect 76894 496848 76899 496904
rect 76116 496846 76899 496848
rect 76116 496844 76122 496846
rect 76833 496843 76899 496846
rect 78438 496844 78444 496908
rect 78508 496906 78514 496908
rect 78581 496906 78647 496909
rect 78508 496904 78647 496906
rect 78508 496848 78586 496904
rect 78642 496848 78647 496904
rect 78508 496846 78647 496848
rect 78508 496844 78514 496846
rect 78581 496843 78647 496846
rect 79174 496844 79180 496908
rect 79244 496906 79250 496908
rect 79409 496906 79475 496909
rect 79244 496904 79475 496906
rect 79244 496848 79414 496904
rect 79470 496848 79475 496904
rect 79244 496846 79475 496848
rect 79244 496844 79250 496846
rect 79409 496843 79475 496846
rect 81014 496844 81020 496908
rect 81084 496906 81090 496908
rect 81341 496906 81407 496909
rect 81084 496904 81407 496906
rect 81084 496848 81346 496904
rect 81402 496848 81407 496904
rect 81084 496846 81407 496848
rect 81084 496844 81090 496846
rect 81341 496843 81407 496846
rect 83590 496844 83596 496908
rect 83660 496906 83666 496908
rect 84101 496906 84167 496909
rect 83660 496904 84167 496906
rect 83660 496848 84106 496904
rect 84162 496848 84167 496904
rect 83660 496846 84167 496848
rect 83660 496844 83666 496846
rect 84101 496843 84167 496846
rect 85982 496844 85988 496908
rect 86052 496906 86058 496908
rect 86861 496906 86927 496909
rect 88241 496908 88307 496909
rect 91001 496908 91067 496909
rect 86052 496904 86927 496906
rect 86052 496848 86866 496904
rect 86922 496848 86927 496904
rect 86052 496846 86927 496848
rect 86052 496844 86058 496846
rect 86861 496843 86927 496846
rect 88190 496844 88196 496908
rect 88260 496906 88307 496908
rect 90950 496906 90956 496908
rect 88260 496904 88352 496906
rect 88302 496848 88352 496904
rect 88260 496846 88352 496848
rect 90910 496846 90956 496906
rect 91020 496904 91067 496908
rect 91062 496848 91067 496904
rect 88260 496844 88307 496846
rect 90950 496844 90956 496846
rect 91020 496844 91067 496848
rect 93526 496844 93532 496908
rect 93596 496906 93602 496908
rect 93761 496906 93827 496909
rect 93596 496904 93827 496906
rect 93596 496848 93766 496904
rect 93822 496848 93827 496904
rect 93596 496846 93827 496848
rect 93596 496844 93602 496846
rect 88241 496843 88307 496844
rect 91001 496843 91067 496844
rect 93761 496843 93827 496846
rect 95918 496844 95924 496908
rect 95988 496906 95994 496908
rect 96521 496906 96587 496909
rect 95988 496904 96587 496906
rect 95988 496848 96526 496904
rect 96582 496848 96587 496904
rect 95988 496846 96587 496848
rect 95988 496844 95994 496846
rect 96521 496843 96587 496846
rect 98494 496844 98500 496908
rect 98564 496906 98570 496908
rect 99281 496906 99347 496909
rect 100937 496908 101003 496909
rect 100886 496906 100892 496908
rect 98564 496904 99347 496906
rect 98564 496848 99286 496904
rect 99342 496848 99347 496904
rect 98564 496846 99347 496848
rect 100846 496846 100892 496906
rect 100956 496904 101003 496908
rect 100998 496848 101003 496904
rect 98564 496844 98570 496846
rect 99281 496843 99347 496846
rect 100886 496844 100892 496846
rect 100956 496844 101003 496848
rect 103462 496844 103468 496908
rect 103532 496906 103538 496908
rect 104801 496906 104867 496909
rect 103532 496904 104867 496906
rect 103532 496848 104806 496904
rect 104862 496848 104867 496904
rect 103532 496846 104867 496848
rect 103532 496844 103538 496846
rect 100937 496843 101003 496844
rect 104801 496843 104867 496846
rect 108614 496844 108620 496908
rect 108684 496906 108690 496908
rect 108849 496906 108915 496909
rect 108684 496904 108915 496906
rect 108684 496848 108854 496904
rect 108910 496848 108915 496904
rect 108684 496846 108915 496848
rect 108684 496844 108690 496846
rect 108849 496843 108915 496846
rect 111006 496844 111012 496908
rect 111076 496906 111082 496908
rect 111701 496906 111767 496909
rect 115841 496908 115907 496909
rect 118601 496908 118667 496909
rect 111076 496904 111767 496906
rect 111076 496848 111706 496904
rect 111762 496848 111767 496904
rect 111076 496846 111767 496848
rect 111076 496844 111082 496846
rect 111701 496843 111767 496846
rect 115790 496844 115796 496908
rect 115860 496906 115907 496908
rect 118550 496906 118556 496908
rect 115860 496904 115952 496906
rect 115902 496848 115952 496904
rect 115860 496846 115952 496848
rect 118510 496846 118556 496906
rect 118620 496904 118667 496908
rect 118662 496848 118667 496904
rect 115860 496844 115907 496846
rect 118550 496844 118556 496846
rect 118620 496844 118667 496848
rect 123334 496844 123340 496908
rect 123404 496906 123410 496908
rect 124121 496906 124187 496909
rect 123404 496904 124187 496906
rect 123404 496848 124126 496904
rect 124182 496848 124187 496904
rect 123404 496846 124187 496848
rect 123404 496844 123410 496846
rect 115841 496843 115907 496844
rect 118601 496843 118667 496844
rect 124121 496843 124187 496846
rect 125910 496844 125916 496908
rect 125980 496906 125986 496908
rect 126881 496906 126947 496909
rect 436093 496908 436159 496909
rect 436093 496906 436140 496908
rect 125980 496904 126947 496906
rect 125980 496848 126886 496904
rect 126942 496848 126947 496904
rect 125980 496846 126947 496848
rect 436048 496904 436140 496906
rect 436048 496848 436098 496904
rect 436048 496846 436140 496848
rect 125980 496844 125986 496846
rect 126881 496843 126947 496846
rect 436093 496844 436140 496846
rect 436204 496844 436210 496908
rect 437473 496906 437539 496909
rect 438342 496906 438348 496908
rect 437473 496904 438348 496906
rect 437473 496848 437478 496904
rect 437534 496848 438348 496904
rect 437473 496846 438348 496848
rect 436093 496843 436159 496844
rect 437473 496843 437539 496846
rect 438342 496844 438348 496846
rect 438412 496844 438418 496908
rect 438853 496906 438919 496909
rect 439630 496906 439636 496908
rect 438853 496904 439636 496906
rect 438853 496848 438858 496904
rect 438914 496848 439636 496904
rect 438853 496846 439636 496848
rect 438853 496843 438919 496846
rect 439630 496844 439636 496846
rect 439700 496844 439706 496908
rect 440233 496906 440299 496909
rect 440550 496906 440556 496908
rect 440233 496904 440556 496906
rect 440233 496848 440238 496904
rect 440294 496848 440556 496904
rect 440233 496846 440556 496848
rect 440233 496843 440299 496846
rect 440550 496844 440556 496846
rect 440620 496844 440626 496908
rect 443126 496844 443132 496908
rect 443196 496906 443202 496908
rect 443637 496906 443703 496909
rect 443196 496904 443703 496906
rect 443196 496848 443642 496904
rect 443698 496848 443703 496904
rect 443196 496846 443703 496848
rect 443196 496844 443202 496846
rect 443637 496843 443703 496846
rect 447133 496906 447199 496909
rect 448278 496906 448284 496908
rect 447133 496904 448284 496906
rect 447133 496848 447138 496904
rect 447194 496848 448284 496904
rect 447133 496846 448284 496848
rect 447133 496843 447199 496846
rect 448278 496844 448284 496846
rect 448348 496844 448354 496908
rect 449893 496906 449959 496909
rect 450670 496906 450676 496908
rect 449893 496904 450676 496906
rect 449893 496848 449898 496904
rect 449954 496848 450676 496904
rect 449893 496846 450676 496848
rect 449893 496843 449959 496846
rect 450670 496844 450676 496846
rect 450740 496844 450746 496908
rect 452653 496906 452719 496909
rect 453614 496906 453620 496908
rect 452653 496904 453620 496906
rect 452653 496848 452658 496904
rect 452714 496848 453620 496904
rect 452653 496846 453620 496848
rect 452653 496843 452719 496846
rect 453614 496844 453620 496846
rect 453684 496844 453690 496908
rect 455822 496844 455828 496908
rect 455892 496906 455898 496908
rect 456057 496906 456123 496909
rect 455892 496904 456123 496906
rect 455892 496848 456062 496904
rect 456118 496848 456123 496904
rect 455892 496846 456123 496848
rect 455892 496844 455898 496846
rect 456057 496843 456123 496846
rect 456885 496908 456994 496909
rect 456885 496904 456932 496908
rect 456996 496906 457002 496908
rect 458173 496906 458239 496909
rect 459461 496908 459527 496909
rect 460933 496908 460999 496909
rect 458398 496906 458404 496908
rect 456885 496848 456890 496904
rect 456885 496844 456932 496848
rect 456996 496846 457042 496906
rect 458173 496904 458404 496906
rect 458173 496848 458178 496904
rect 458234 496848 458404 496904
rect 458173 496846 458404 496848
rect 456996 496844 457002 496846
rect 456885 496843 456951 496844
rect 458173 496843 458239 496846
rect 458398 496844 458404 496846
rect 458468 496844 458474 496908
rect 459461 496904 459508 496908
rect 459572 496906 459578 496908
rect 459461 496848 459466 496904
rect 459461 496844 459508 496848
rect 459572 496846 459618 496906
rect 460933 496904 460980 496908
rect 461044 496906 461050 496908
rect 462405 496906 462471 496909
rect 463550 496906 463556 496908
rect 460933 496848 460938 496904
rect 459572 496844 459578 496846
rect 460933 496844 460980 496848
rect 461044 496846 461090 496906
rect 462405 496904 463556 496906
rect 462405 496848 462410 496904
rect 462466 496848 463556 496904
rect 462405 496846 463556 496848
rect 461044 496844 461050 496846
rect 459461 496843 459527 496844
rect 460933 496843 460999 496844
rect 462405 496843 462471 496846
rect 463550 496844 463556 496846
rect 463620 496844 463626 496908
rect 465165 496906 465231 496909
rect 465942 496906 465948 496908
rect 465165 496904 465948 496906
rect 465165 496848 465170 496904
rect 465226 496848 465948 496904
rect 465165 496846 465948 496848
rect 465165 496843 465231 496846
rect 465942 496844 465948 496846
rect 466012 496844 466018 496908
rect 467925 496906 467991 496909
rect 468334 496906 468340 496908
rect 467925 496904 468340 496906
rect 467925 496848 467930 496904
rect 467986 496848 468340 496904
rect 467925 496846 468340 496848
rect 467925 496843 467991 496846
rect 468334 496844 468340 496846
rect 468404 496844 468410 496908
rect 470777 496906 470843 496909
rect 476113 496908 476179 496909
rect 470910 496906 470916 496908
rect 470777 496904 470916 496906
rect 470777 496848 470782 496904
rect 470838 496848 470916 496904
rect 470777 496846 470916 496848
rect 470777 496843 470843 496846
rect 470910 496844 470916 496846
rect 470980 496844 470986 496908
rect 476062 496906 476068 496908
rect 476022 496846 476068 496906
rect 476132 496904 476179 496908
rect 476174 496848 476179 496904
rect 476062 496844 476068 496846
rect 476132 496844 476179 496848
rect 476113 496843 476179 496844
rect 477493 496906 477559 496909
rect 478086 496906 478092 496908
rect 477493 496904 478092 496906
rect 477493 496848 477498 496904
rect 477554 496848 478092 496904
rect 477493 496846 478092 496848
rect 477493 496843 477559 496846
rect 478086 496844 478092 496846
rect 478156 496844 478162 496908
rect 483013 496906 483079 496909
rect 483422 496906 483428 496908
rect 483013 496904 483428 496906
rect 483013 496848 483018 496904
rect 483074 496848 483428 496904
rect 483013 496846 483428 496848
rect 483013 496843 483079 496846
rect 483422 496844 483428 496846
rect 483492 496844 483498 496908
rect 485773 496906 485839 496909
rect 485998 496906 486004 496908
rect 485773 496904 486004 496906
rect 485773 496848 485778 496904
rect 485834 496848 486004 496904
rect 485773 496846 486004 496848
rect 485773 496843 485839 496846
rect 485998 496844 486004 496846
rect 486068 496844 486074 496908
rect 487153 496906 487219 496909
rect 488206 496906 488212 496908
rect 487153 496904 488212 496906
rect 487153 496848 487158 496904
rect 487214 496848 488212 496904
rect 487153 496846 488212 496848
rect 487153 496843 487219 496846
rect 488206 496844 488212 496846
rect 488276 496844 488282 496908
rect 490465 496906 490531 496909
rect 490966 496906 490972 496908
rect 490465 496904 490972 496906
rect 490465 496848 490470 496904
rect 490526 496848 490972 496904
rect 490465 496846 490972 496848
rect 490465 496843 490531 496846
rect 490966 496844 490972 496846
rect 491036 496844 491042 496908
rect 492673 496906 492739 496909
rect 493358 496906 493364 496908
rect 492673 496904 493364 496906
rect 492673 496848 492678 496904
rect 492734 496848 493364 496904
rect 492673 496846 493364 496848
rect 492673 496843 492739 496846
rect 493358 496844 493364 496846
rect 493428 496844 493434 496908
rect 497457 496906 497523 496909
rect 500953 496908 501019 496909
rect 498510 496906 498516 496908
rect 497457 496904 498516 496906
rect 497457 496848 497462 496904
rect 497518 496848 498516 496904
rect 497457 496846 498516 496848
rect 497457 496843 497523 496846
rect 498510 496844 498516 496846
rect 498580 496844 498586 496908
rect 500902 496906 500908 496908
rect 500862 496846 500908 496906
rect 500972 496904 501019 496908
rect 501014 496848 501019 496904
rect 500902 496844 500908 496846
rect 500972 496844 501019 496848
rect 500953 496843 501019 496844
rect 502333 496906 502399 496909
rect 503478 496906 503484 496908
rect 502333 496904 503484 496906
rect 502333 496848 502338 496904
rect 502394 496848 503484 496904
rect 502333 496846 503484 496848
rect 502333 496843 502399 496846
rect 503478 496844 503484 496846
rect 503548 496844 503554 496908
rect 507853 496906 507919 496909
rect 508446 496906 508452 496908
rect 507853 496904 508452 496906
rect 507853 496848 507858 496904
rect 507914 496848 508452 496904
rect 507853 496846 508452 496848
rect 507853 496843 507919 496846
rect 508446 496844 508452 496846
rect 508516 496844 508522 496908
rect 510613 496906 510679 496909
rect 511022 496906 511028 496908
rect 510613 496904 511028 496906
rect 510613 496848 510618 496904
rect 510674 496848 511028 496904
rect 510613 496846 511028 496848
rect 510613 496843 510679 496846
rect 511022 496844 511028 496846
rect 511092 496844 511098 496908
rect 514753 496906 514819 496909
rect 515806 496906 515812 496908
rect 514753 496904 515812 496906
rect 514753 496848 514758 496904
rect 514814 496848 515812 496904
rect 514753 496846 515812 496848
rect 514753 496843 514819 496846
rect 515806 496844 515812 496846
rect 515876 496844 515882 496908
rect 517513 496906 517579 496909
rect 518382 496906 518388 496908
rect 517513 496904 518388 496906
rect 517513 496848 517518 496904
rect 517574 496848 518388 496904
rect 517513 496846 518388 496848
rect 517513 496843 517579 496846
rect 518382 496844 518388 496846
rect 518452 496844 518458 496908
rect 523033 496906 523099 496909
rect 523350 496906 523356 496908
rect 523033 496904 523356 496906
rect 523033 496848 523038 496904
rect 523094 496848 523356 496904
rect 523033 496846 523356 496848
rect 523033 496843 523099 496846
rect 523350 496844 523356 496846
rect 523420 496844 523426 496908
rect 525793 496906 525859 496909
rect 525926 496906 525932 496908
rect 525793 496904 525932 496906
rect 525793 496848 525798 496904
rect 525854 496848 525932 496904
rect 525793 496846 525932 496848
rect 525793 496843 525859 496846
rect 525926 496844 525932 496846
rect 525996 496844 526002 496908
rect 418705 496770 418771 496773
rect 419758 496770 419764 496772
rect 418705 496768 419764 496770
rect 418705 496712 418710 496768
rect 418766 496712 419764 496768
rect 418705 496710 419764 496712
rect 418705 496707 418771 496710
rect 419758 496708 419764 496710
rect 419828 496770 419834 496772
rect 420729 496770 420795 496773
rect 419828 496768 420795 496770
rect 419828 496712 420734 496768
rect 420790 496712 420795 496768
rect 419828 496710 420795 496712
rect 419828 496708 419834 496710
rect 420729 496707 420795 496710
rect 18638 496028 18644 496092
rect 18708 496090 18714 496092
rect 277393 496090 277459 496093
rect 18708 496088 277459 496090
rect 18708 496032 277398 496088
rect 277454 496032 277459 496088
rect 18708 496030 277459 496032
rect 18708 496028 18714 496030
rect 277393 496027 277459 496030
rect 259729 495002 259795 495005
rect 374126 495002 374132 495004
rect 259729 495000 374132 495002
rect 259729 494944 259734 495000
rect 259790 494944 374132 495000
rect 259729 494942 374132 494944
rect 259729 494939 259795 494942
rect 374126 494940 374132 494942
rect 374196 494940 374202 495004
rect 244457 494866 244523 494869
rect 372654 494866 372660 494868
rect 244457 494864 372660 494866
rect 244457 494808 244462 494864
rect 244518 494808 372660 494864
rect 244457 494806 372660 494808
rect 244457 494803 244523 494806
rect 372654 494804 372660 494806
rect 372724 494804 372730 494868
rect 19006 494668 19012 494732
rect 19076 494730 19082 494732
rect 41873 494730 41939 494733
rect 19076 494728 41939 494730
rect 19076 494672 41878 494728
rect 41934 494672 41939 494728
rect 19076 494670 41939 494672
rect 19076 494668 19082 494670
rect 41873 494667 41939 494670
rect 245745 494730 245811 494733
rect 373758 494730 373764 494732
rect 245745 494728 373764 494730
rect 245745 494672 245750 494728
rect 245806 494672 373764 494728
rect 245745 494670 373764 494672
rect 245745 494667 245811 494670
rect 373758 494668 373764 494670
rect 373828 494668 373834 494732
rect 416681 494050 416747 494053
rect 417366 494050 417372 494052
rect 416681 494048 417372 494050
rect 416681 493992 416686 494048
rect 416742 493992 417372 494048
rect 416681 493990 417372 493992
rect 416681 493987 416747 493990
rect 417366 493988 417372 493990
rect 417436 494050 417442 494052
rect 441613 494050 441679 494053
rect 417436 494048 441679 494050
rect 417436 493992 441618 494048
rect 441674 493992 441679 494048
rect 417436 493990 441679 493992
rect 417436 493988 417442 493990
rect 441613 493987 441679 493990
rect 280153 493370 280219 493373
rect 418838 493370 418844 493372
rect 280153 493368 418844 493370
rect 280153 493312 280158 493368
rect 280214 493312 418844 493368
rect 280153 493310 418844 493312
rect 280153 493307 280219 493310
rect 418838 493308 418844 493310
rect 418908 493308 418914 493372
rect 19149 491194 19215 491197
rect 19742 491194 19748 491196
rect 19149 491192 19748 491194
rect 19149 491136 19154 491192
rect 19210 491136 19748 491192
rect 19149 491134 19748 491136
rect 19149 491131 19215 491134
rect 19742 491132 19748 491134
rect 19812 491194 19818 491196
rect 37273 491194 37339 491197
rect 19812 491192 37339 491194
rect 19812 491136 37278 491192
rect 37334 491136 37339 491192
rect 19812 491134 37339 491136
rect 19812 491132 19818 491134
rect 37273 491131 37339 491134
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 209865 480858 209931 480861
rect 418654 480858 418660 480860
rect 209865 480856 418660 480858
rect 209865 480800 209870 480856
rect 209926 480800 418660 480856
rect 209865 480798 418660 480800
rect 209865 480795 209931 480798
rect 418654 480796 418660 480798
rect 418724 480796 418730 480860
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 195094 475356 195100 475420
rect 195164 475418 195170 475420
rect 338205 475418 338271 475421
rect 195164 475416 338271 475418
rect 195164 475360 338210 475416
rect 338266 475360 338271 475416
rect 195164 475358 338271 475360
rect 195164 475356 195170 475358
rect 338205 475355 338271 475358
rect 15929 474058 15995 474061
rect 287697 474058 287763 474061
rect 15929 474056 287763 474058
rect 15929 474000 15934 474056
rect 15990 474000 287702 474056
rect 287758 474000 287763 474056
rect 15929 473998 287763 474000
rect 15929 473995 15995 473998
rect 287697 473995 287763 473998
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 199326 468420 199332 468484
rect 199396 468482 199402 468484
rect 218053 468482 218119 468485
rect 199396 468480 218119 468482
rect 199396 468424 218058 468480
rect 218114 468424 218119 468480
rect 199396 468422 218119 468424
rect 199396 468420 199402 468422
rect 218053 468419 218119 468422
rect 203558 466108 203564 466172
rect 203628 466170 203634 466172
rect 248597 466170 248663 466173
rect 203628 466168 248663 466170
rect 203628 466112 248602 466168
rect 248658 466112 248663 466168
rect 203628 466110 248663 466112
rect 203628 466108 203634 466110
rect 248597 466107 248663 466110
rect 197813 466034 197879 466037
rect 314653 466034 314719 466037
rect 197813 466032 314719 466034
rect 197813 465976 197818 466032
rect 197874 465976 314658 466032
rect 314714 465976 314719 466032
rect 197813 465974 314719 465976
rect 197813 465971 197879 465974
rect 314653 465971 314719 465974
rect 198038 465836 198044 465900
rect 198108 465898 198114 465900
rect 317413 465898 317479 465901
rect 198108 465896 317479 465898
rect 198108 465840 317418 465896
rect 317474 465840 317479 465896
rect 198108 465838 317479 465840
rect 198108 465836 198114 465838
rect 317413 465835 317479 465838
rect 156689 465762 156755 465765
rect 385125 465762 385191 465765
rect 156689 465760 385191 465762
rect 156689 465704 156694 465760
rect 156750 465704 385130 465760
rect 385186 465704 385191 465760
rect 156689 465702 385191 465704
rect 156689 465699 156755 465702
rect 385125 465699 385191 465702
rect 192702 463660 192708 463724
rect 192772 463722 192778 463724
rect 273253 463722 273319 463725
rect 417417 463724 417483 463725
rect 417366 463722 417372 463724
rect 192772 463720 273319 463722
rect 192772 463664 273258 463720
rect 273314 463664 273319 463720
rect 192772 463662 273319 463664
rect 417326 463662 417372 463722
rect 417436 463720 417483 463724
rect 417478 463664 417483 463720
rect 192772 463660 192778 463662
rect 273253 463659 273319 463662
rect 417366 463660 417372 463662
rect 417436 463660 417483 463664
rect 417417 463659 417483 463660
rect 173341 463042 173407 463045
rect 302325 463042 302391 463045
rect 173341 463040 302391 463042
rect 173341 462984 173346 463040
rect 173402 462984 302330 463040
rect 302386 462984 302391 463040
rect 173341 462982 302391 462984
rect 173341 462979 173407 462982
rect 302325 462979 302391 462982
rect 211337 462906 211403 462909
rect 393957 462906 394023 462909
rect 211337 462904 394023 462906
rect 211337 462848 211342 462904
rect 211398 462848 393962 462904
rect 394018 462848 394023 462904
rect 211337 462846 394023 462848
rect 211337 462843 211403 462846
rect 393957 462843 394023 462846
rect 173157 462770 173223 462773
rect 310697 462770 310763 462773
rect 173157 462768 310763 462770
rect -960 462634 480 462724
rect 173157 462712 173162 462768
rect 173218 462712 310702 462768
rect 310758 462712 310763 462768
rect 173157 462710 310763 462712
rect 173157 462707 173223 462710
rect 310697 462707 310763 462710
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 170397 462634 170463 462637
rect 317505 462634 317571 462637
rect 170397 462632 317571 462634
rect 170397 462576 170402 462632
rect 170458 462576 317510 462632
rect 317566 462576 317571 462632
rect 170397 462574 317571 462576
rect 170397 462571 170463 462574
rect 317505 462571 317571 462574
rect 175917 462498 175983 462501
rect 364425 462498 364491 462501
rect 175917 462496 364491 462498
rect 175917 462440 175922 462496
rect 175978 462440 364430 462496
rect 364486 462440 364491 462496
rect 175917 462438 364491 462440
rect 175917 462435 175983 462438
rect 364425 462435 364491 462438
rect 173525 462362 173591 462365
rect 379605 462362 379671 462365
rect 173525 462360 379671 462362
rect 173525 462304 173530 462360
rect 173586 462304 379610 462360
rect 379666 462304 379671 462360
rect 173525 462302 379671 462304
rect 173525 462299 173591 462302
rect 379605 462299 379671 462302
rect 199878 461620 199884 461684
rect 199948 461682 199954 461684
rect 376845 461682 376911 461685
rect 199948 461680 376911 461682
rect 199948 461624 376850 461680
rect 376906 461624 376911 461680
rect 199948 461622 376911 461624
rect 199948 461620 199954 461622
rect 376845 461619 376911 461622
rect 201350 461484 201356 461548
rect 201420 461546 201426 461548
rect 379697 461546 379763 461549
rect 201420 461544 379763 461546
rect 201420 461488 379702 461544
rect 379758 461488 379763 461544
rect 201420 461486 379763 461488
rect 201420 461484 201426 461486
rect 379697 461483 379763 461486
rect 192150 461348 192156 461412
rect 192220 461410 192226 461412
rect 272149 461410 272215 461413
rect 192220 461408 272215 461410
rect 192220 461352 272154 461408
rect 272210 461352 272215 461408
rect 192220 461350 272215 461352
rect 192220 461348 192226 461350
rect 272149 461347 272215 461350
rect 173249 461274 173315 461277
rect 314745 461274 314811 461277
rect 173249 461272 314811 461274
rect 173249 461216 173254 461272
rect 173310 461216 314750 461272
rect 314806 461216 314811 461272
rect 173249 461214 314811 461216
rect 173249 461211 173315 461214
rect 314745 461211 314811 461214
rect 176101 461138 176167 461141
rect 370129 461138 370195 461141
rect 176101 461136 370195 461138
rect 176101 461080 176106 461136
rect 176162 461080 370134 461136
rect 370190 461080 370195 461136
rect 176101 461078 370195 461080
rect 176101 461075 176167 461078
rect 370129 461075 370195 461078
rect 173709 461002 173775 461005
rect 375465 461002 375531 461005
rect 173709 461000 375531 461002
rect 173709 460944 173714 461000
rect 173770 460944 375470 461000
rect 375526 460944 375531 461000
rect 173709 460942 375531 460944
rect 173709 460939 173775 460942
rect 375465 460939 375531 460942
rect 179321 460322 179387 460325
rect 331397 460322 331463 460325
rect 179321 460320 331463 460322
rect 179321 460264 179326 460320
rect 179382 460264 331402 460320
rect 331458 460264 331463 460320
rect 179321 460262 331463 460264
rect 179321 460259 179387 460262
rect 331397 460259 331463 460262
rect 197854 460124 197860 460188
rect 197924 460186 197930 460188
rect 382549 460186 382615 460189
rect 197924 460184 382615 460186
rect 197924 460128 382554 460184
rect 382610 460128 382615 460184
rect 197924 460126 382615 460128
rect 197924 460124 197930 460126
rect 382549 460123 382615 460126
rect 179137 460050 179203 460053
rect 337653 460050 337719 460053
rect 179137 460048 337719 460050
rect 179137 459992 179142 460048
rect 179198 459992 337658 460048
rect 337714 459992 337719 460048
rect 179137 459990 337719 459992
rect 179137 459987 179203 459990
rect 337653 459987 337719 459990
rect 178585 459914 178651 459917
rect 343909 459914 343975 459917
rect 178585 459912 343975 459914
rect 178585 459856 178590 459912
rect 178646 459856 343914 459912
rect 343970 459856 343975 459912
rect 178585 459854 343975 459856
rect 178585 459851 178651 459854
rect 343909 459851 343975 459854
rect 176009 459778 176075 459781
rect 352741 459778 352807 459781
rect 176009 459776 352807 459778
rect 176009 459720 176014 459776
rect 176070 459720 352746 459776
rect 352802 459720 352807 459776
rect 176009 459718 352807 459720
rect 176009 459715 176075 459718
rect 352741 459715 352807 459718
rect 176193 459642 176259 459645
rect 358997 459642 359063 459645
rect 176193 459640 359063 459642
rect 176193 459584 176198 459640
rect 176254 459584 359002 459640
rect 359058 459584 359063 459640
rect 176193 459582 359063 459584
rect 176193 459579 176259 459582
rect 358997 459579 359063 459582
rect 188470 458900 188476 458964
rect 188540 458962 188546 458964
rect 309317 458962 309383 458965
rect 188540 458960 309383 458962
rect 188540 458904 309322 458960
rect 309378 458904 309383 458960
rect 188540 458902 309383 458904
rect 188540 458900 188546 458902
rect 309317 458899 309383 458902
rect 178953 458826 179019 458829
rect 346853 458826 346919 458829
rect 178953 458824 346919 458826
rect 178953 458768 178958 458824
rect 179014 458768 346858 458824
rect 346914 458768 346919 458824
rect 178953 458766 346919 458768
rect 178953 458763 179019 458766
rect 346853 458763 346919 458766
rect 176285 458690 176351 458693
rect 355685 458690 355751 458693
rect 176285 458688 355751 458690
rect 176285 458632 176290 458688
rect 176346 458632 355690 458688
rect 355746 458632 355751 458688
rect 176285 458630 355751 458632
rect 176285 458627 176351 458630
rect 355685 458627 355751 458630
rect 176469 458554 176535 458557
rect 361665 458554 361731 458557
rect 176469 458552 361731 458554
rect 176469 458496 176474 458552
rect 176530 458496 361670 458552
rect 361726 458496 361731 458552
rect 176469 458494 361731 458496
rect 176469 458491 176535 458494
rect 361665 458491 361731 458494
rect 197537 458418 197603 458421
rect 580533 458418 580599 458421
rect 197537 458416 580599 458418
rect 197537 458360 197542 458416
rect 197598 458360 580538 458416
rect 580594 458360 580599 458416
rect 197537 458358 580599 458360
rect 197537 458355 197603 458358
rect 580533 458355 580599 458358
rect 195973 458282 196039 458285
rect 580349 458282 580415 458285
rect 195973 458280 580415 458282
rect 195973 458224 195978 458280
rect 196034 458224 580354 458280
rect 580410 458224 580415 458280
rect 195973 458222 580415 458224
rect 195973 458219 196039 458222
rect 580349 458219 580415 458222
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 176377 457602 176443 457605
rect 285949 457602 286015 457605
rect 176377 457600 286015 457602
rect 176377 457544 176382 457600
rect 176438 457544 285954 457600
rect 286010 457544 286015 457600
rect 176377 457542 286015 457544
rect 176377 457539 176443 457542
rect 285949 457539 286015 457542
rect 211429 457466 211495 457469
rect 415894 457466 415900 457468
rect 211429 457464 415900 457466
rect 211429 457408 211434 457464
rect 211490 457408 415900 457464
rect 211429 457406 415900 457408
rect 211429 457403 211495 457406
rect 415894 457404 415900 457406
rect 415964 457404 415970 457468
rect 186814 457268 186820 457332
rect 186884 457330 186890 457332
rect 342529 457330 342595 457333
rect 186884 457328 342595 457330
rect 186884 457272 342534 457328
rect 342590 457272 342595 457328
rect 186884 457270 342595 457272
rect 186884 457268 186890 457270
rect 342529 457267 342595 457270
rect 184054 457132 184060 457196
rect 184124 457194 184130 457196
rect 371877 457194 371943 457197
rect 184124 457192 371943 457194
rect 184124 457136 371882 457192
rect 371938 457136 371943 457192
rect 184124 457134 371943 457136
rect 184124 457132 184130 457134
rect 371877 457131 371943 457134
rect 181805 457058 181871 457061
rect 377765 457058 377831 457061
rect 181805 457056 377831 457058
rect 181805 457000 181810 457056
rect 181866 457000 377770 457056
rect 377826 457000 377831 457056
rect 181805 456998 377831 457000
rect 181805 456995 181871 456998
rect 377765 456995 377831 456998
rect 19190 456860 19196 456924
rect 19260 456922 19266 456924
rect 283005 456922 283071 456925
rect 19260 456920 283071 456922
rect 19260 456864 283010 456920
rect 283066 456864 283071 456920
rect 19260 456862 283071 456864
rect 19260 456860 19266 456862
rect 283005 456859 283071 456862
rect 173801 456242 173867 456245
rect 289997 456242 290063 456245
rect 173801 456240 290063 456242
rect 173801 456184 173806 456240
rect 173862 456184 290002 456240
rect 290058 456184 290063 456240
rect 173801 456182 290063 456184
rect 173801 456179 173867 456182
rect 289997 456179 290063 456182
rect 186998 456044 187004 456108
rect 187068 456106 187074 456108
rect 332869 456106 332935 456109
rect 187068 456104 332935 456106
rect 187068 456048 332874 456104
rect 332930 456048 332935 456104
rect 187068 456046 332935 456048
rect 187068 456044 187074 456046
rect 332869 456043 332935 456046
rect 187182 455908 187188 455972
rect 187252 455970 187258 455972
rect 348325 455970 348391 455973
rect 187252 455968 348391 455970
rect 187252 455912 348330 455968
rect 348386 455912 348391 455968
rect 187252 455910 348391 455912
rect 187252 455908 187258 455910
rect 348325 455907 348391 455910
rect 184238 455772 184244 455836
rect 184308 455834 184314 455836
rect 375097 455834 375163 455837
rect 184308 455832 375163 455834
rect 184308 455776 375102 455832
rect 375158 455776 375163 455832
rect 184308 455774 375163 455776
rect 184308 455772 184314 455774
rect 375097 455771 375163 455774
rect 197353 455698 197419 455701
rect 573357 455698 573423 455701
rect 197353 455696 573423 455698
rect 197353 455640 197358 455696
rect 197414 455640 573362 455696
rect 573418 455640 573423 455696
rect 197353 455638 573423 455640
rect 197353 455635 197419 455638
rect 573357 455635 573423 455638
rect 196249 455562 196315 455565
rect 571977 455562 572043 455565
rect 196249 455560 572043 455562
rect 196249 455504 196254 455560
rect 196310 455504 571982 455560
rect 572038 455504 572043 455560
rect 196249 455502 572043 455504
rect 196249 455499 196315 455502
rect 571977 455499 572043 455502
rect 190310 454684 190316 454748
rect 190380 454746 190386 454748
rect 277669 454746 277735 454749
rect 190380 454744 277735 454746
rect 190380 454688 277674 454744
rect 277730 454688 277735 454744
rect 190380 454686 277735 454688
rect 190380 454684 190386 454686
rect 277669 454683 277735 454686
rect 188286 454548 188292 454612
rect 188356 454610 188362 454612
rect 373625 454610 373691 454613
rect 188356 454608 373691 454610
rect 188356 454552 373630 454608
rect 373686 454552 373691 454608
rect 188356 454550 373691 454552
rect 188356 454548 188362 454550
rect 373625 454547 373691 454550
rect 191046 454412 191052 454476
rect 191116 454474 191122 454476
rect 382365 454474 382431 454477
rect 191116 454472 382431 454474
rect 191116 454416 382370 454472
rect 382426 454416 382431 454472
rect 191116 454414 382431 454416
rect 191116 454412 191122 454414
rect 382365 454411 382431 454414
rect 18454 454276 18460 454340
rect 18524 454338 18530 454340
rect 232773 454338 232839 454341
rect 18524 454336 232839 454338
rect 18524 454280 232778 454336
rect 232834 454280 232839 454336
rect 18524 454278 232839 454280
rect 18524 454276 18530 454278
rect 232773 454275 232839 454278
rect 289077 454338 289143 454341
rect 414606 454338 414612 454340
rect 289077 454336 414612 454338
rect 289077 454280 289082 454336
rect 289138 454280 414612 454336
rect 289077 454278 414612 454280
rect 289077 454275 289143 454278
rect 414606 454276 414612 454278
rect 414676 454276 414682 454340
rect 194593 454202 194659 454205
rect 558177 454202 558243 454205
rect 194593 454200 558243 454202
rect 194593 454144 194598 454200
rect 194654 454144 558182 454200
rect 558238 454144 558243 454200
rect 194593 454142 558243 454144
rect 194593 454139 194659 454142
rect 558177 454139 558243 454142
rect 196985 454066 197051 454069
rect 566457 454066 566523 454069
rect 196985 454064 566523 454066
rect 196985 454008 196990 454064
rect 197046 454008 566462 454064
rect 566518 454008 566523 454064
rect 196985 454006 566523 454008
rect 196985 454003 197051 454006
rect 566457 454003 566523 454006
rect 187325 453386 187391 453389
rect 230105 453386 230171 453389
rect 187325 453384 230171 453386
rect 187325 453328 187330 453384
rect 187386 453328 230110 453384
rect 230166 453328 230171 453384
rect 187325 453326 230171 453328
rect 187325 453323 187391 453326
rect 230105 453323 230171 453326
rect 185158 453188 185164 453252
rect 185228 453250 185234 453252
rect 265433 453250 265499 453253
rect 185228 453248 265499 453250
rect 185228 453192 265438 453248
rect 265494 453192 265499 453248
rect 185228 453190 265499 453192
rect 185228 453188 185234 453190
rect 265433 453187 265499 453190
rect 192518 453052 192524 453116
rect 192588 453114 192594 453116
rect 273897 453114 273963 453117
rect 192588 453112 273963 453114
rect 192588 453056 273902 453112
rect 273958 453056 273963 453112
rect 192588 453054 273963 453056
rect 192588 453052 192594 453054
rect 273897 453051 273963 453054
rect 284937 453114 285003 453117
rect 418102 453114 418108 453116
rect 284937 453112 418108 453114
rect 284937 453056 284942 453112
rect 284998 453056 418108 453112
rect 284937 453054 418108 453056
rect 284937 453051 285003 453054
rect 418102 453052 418108 453054
rect 418172 453052 418178 453116
rect 176561 452978 176627 452981
rect 350073 452978 350139 452981
rect 176561 452976 350139 452978
rect 176561 452920 176566 452976
rect 176622 452920 350078 452976
rect 350134 452920 350139 452976
rect 176561 452918 350139 452920
rect 176561 452915 176627 452918
rect 350073 452915 350139 452918
rect 18781 452842 18847 452845
rect 300393 452842 300459 452845
rect 18781 452840 300459 452842
rect 18781 452784 18786 452840
rect 18842 452784 300398 452840
rect 300454 452784 300459 452840
rect 18781 452782 300459 452784
rect 18781 452779 18847 452782
rect 300393 452779 300459 452782
rect 193673 452706 193739 452709
rect 580257 452706 580323 452709
rect 193673 452704 580323 452706
rect 193673 452648 193678 452704
rect 193734 452648 580262 452704
rect 580318 452648 580323 452704
rect 193673 452646 580323 452648
rect 193673 452643 193739 452646
rect 580257 452643 580323 452646
rect 248454 452508 248460 452572
rect 248524 452570 248530 452572
rect 248873 452570 248939 452573
rect 248524 452568 248939 452570
rect 248524 452512 248878 452568
rect 248934 452512 248939 452568
rect 248524 452510 248939 452512
rect 248524 452508 248530 452510
rect 248873 452507 248939 452510
rect 373257 452570 373323 452573
rect 374494 452570 374500 452572
rect 373257 452568 374500 452570
rect 373257 452512 373262 452568
rect 373318 452512 374500 452568
rect 373257 452510 374500 452512
rect 373257 452507 373323 452510
rect 374494 452508 374500 452510
rect 374564 452508 374570 452572
rect 376201 452570 376267 452573
rect 376334 452570 376340 452572
rect 376201 452568 376340 452570
rect 376201 452512 376206 452568
rect 376262 452512 376340 452568
rect 376201 452510 376340 452512
rect 376201 452507 376267 452510
rect 376334 452508 376340 452510
rect 376404 452508 376410 452572
rect 369945 452434 370011 452437
rect 418654 452434 418660 452436
rect 369945 452432 418660 452434
rect 369945 452376 369950 452432
rect 370006 452376 418660 452432
rect 369945 452374 418660 452376
rect 369945 452371 370011 452374
rect 418654 452372 418660 452374
rect 418724 452372 418730 452436
rect 3417 452298 3483 452301
rect 234889 452298 234955 452301
rect 3417 452296 234955 452298
rect 3417 452240 3422 452296
rect 3478 452240 234894 452296
rect 234950 452240 234955 452296
rect 3417 452238 234955 452240
rect 3417 452235 3483 452238
rect 234889 452235 234955 452238
rect 375833 452298 375899 452301
rect 418838 452298 418844 452300
rect 375833 452296 418844 452298
rect 375833 452240 375838 452296
rect 375894 452240 418844 452296
rect 375833 452238 418844 452240
rect 375833 452235 375899 452238
rect 418838 452236 418844 452238
rect 418908 452236 418914 452300
rect 203742 452100 203748 452164
rect 203812 452162 203818 452164
rect 235993 452162 236059 452165
rect 203812 452160 236059 452162
rect 203812 452104 235998 452160
rect 236054 452104 236059 452160
rect 203812 452102 236059 452104
rect 203812 452100 203818 452102
rect 235993 452099 236059 452102
rect 364057 452162 364123 452165
rect 368749 452162 368815 452165
rect 364057 452160 368815 452162
rect 364057 452104 364062 452160
rect 364118 452104 368754 452160
rect 368810 452104 368815 452160
rect 364057 452102 368815 452104
rect 364057 452099 364123 452102
rect 368749 452099 368815 452102
rect 190085 452026 190151 452029
rect 264697 452026 264763 452029
rect 190085 452024 264763 452026
rect 190085 451968 190090 452024
rect 190146 451968 264702 452024
rect 264758 451968 264763 452024
rect 190085 451966 264763 451968
rect 190085 451963 190151 451966
rect 264697 451963 264763 451966
rect 352281 452026 352347 452029
rect 378133 452026 378199 452029
rect 352281 452024 378199 452026
rect 352281 451968 352286 452024
rect 352342 451968 378138 452024
rect 378194 451968 378199 452024
rect 352281 451966 378199 451968
rect 352281 451963 352347 451966
rect 378133 451963 378199 451966
rect 189993 451890 190059 451893
rect 266169 451890 266235 451893
rect 189993 451888 266235 451890
rect 189993 451832 189998 451888
rect 190054 451832 266174 451888
rect 266230 451832 266235 451888
rect 189993 451830 266235 451832
rect 189993 451827 190059 451830
rect 266169 451827 266235 451830
rect 300761 451890 300827 451893
rect 372429 451890 372495 451893
rect 300761 451888 372495 451890
rect 300761 451832 300766 451888
rect 300822 451832 372434 451888
rect 372490 451832 372495 451888
rect 300761 451830 372495 451832
rect 300761 451827 300827 451830
rect 372429 451827 372495 451830
rect 378777 451890 378843 451893
rect 415894 451890 415900 451892
rect 378777 451888 415900 451890
rect 378777 451832 378782 451888
rect 378838 451832 415900 451888
rect 378777 451830 415900 451832
rect 378777 451827 378843 451830
rect 415894 451828 415900 451830
rect 415964 451828 415970 451892
rect 188337 451754 188403 451757
rect 266905 451754 266971 451757
rect 188337 451752 266971 451754
rect 188337 451696 188342 451752
rect 188398 451696 266910 451752
rect 266966 451696 266971 451752
rect 188337 451694 266971 451696
rect 188337 451691 188403 451694
rect 266905 451691 266971 451694
rect 319161 451754 319227 451757
rect 419022 451754 419028 451756
rect 319161 451752 419028 451754
rect 319161 451696 319166 451752
rect 319222 451696 419028 451752
rect 319161 451694 419028 451696
rect 319161 451691 319227 451694
rect 419022 451692 419028 451694
rect 419092 451692 419098 451756
rect 184565 451618 184631 451621
rect 284201 451618 284267 451621
rect 184565 451616 284267 451618
rect 184565 451560 184570 451616
rect 184626 451560 284206 451616
rect 284262 451560 284267 451616
rect 184565 451558 284267 451560
rect 184565 451555 184631 451558
rect 284201 451555 284267 451558
rect 292297 451618 292363 451621
rect 408033 451618 408099 451621
rect 292297 451616 408099 451618
rect 292297 451560 292302 451616
rect 292358 451560 408038 451616
rect 408094 451560 408099 451616
rect 292297 451558 408099 451560
rect 292297 451555 292363 451558
rect 408033 451555 408099 451558
rect 188889 451484 188955 451485
rect 188838 451482 188844 451484
rect 188798 451422 188844 451482
rect 188908 451480 188955 451484
rect 195145 451482 195211 451485
rect 188950 451424 188955 451480
rect 188838 451420 188844 451422
rect 188908 451420 188955 451424
rect 188889 451419 188955 451420
rect 190410 451480 195211 451482
rect 190410 451424 195150 451480
rect 195206 451424 195211 451480
rect 190410 451422 195211 451424
rect 188654 451284 188660 451348
rect 188724 451346 188730 451348
rect 190410 451346 190470 451422
rect 195145 451419 195211 451422
rect 201401 451482 201467 451485
rect 390369 451482 390435 451485
rect 201401 451480 390435 451482
rect 201401 451424 201406 451480
rect 201462 451424 390374 451480
rect 390430 451424 390435 451480
rect 201401 451422 390435 451424
rect 201401 451419 201467 451422
rect 390369 451419 390435 451422
rect 188724 451286 190470 451346
rect 188724 451284 188730 451286
rect 191598 451284 191604 451348
rect 191668 451346 191674 451348
rect 195881 451346 195947 451349
rect 191668 451344 195947 451346
rect 191668 451288 195886 451344
rect 195942 451288 195947 451344
rect 191668 451286 195947 451288
rect 191668 451284 191674 451286
rect 195881 451283 195947 451286
rect 287881 451346 287947 451349
rect 410609 451346 410675 451349
rect 287881 451344 410675 451346
rect 287881 451288 287886 451344
rect 287942 451288 410614 451344
rect 410670 451288 410675 451344
rect 287881 451286 410675 451288
rect 287881 451283 287947 451286
rect 410609 451283 410675 451286
rect 383653 450938 383719 450941
rect 417734 450938 417740 450940
rect 383653 450936 417740 450938
rect 383653 450880 383658 450936
rect 383714 450880 417740 450936
rect 383653 450878 417740 450880
rect 383653 450875 383719 450878
rect 417734 450876 417740 450878
rect 417804 450876 417810 450940
rect 191230 450740 191236 450804
rect 191300 450802 191306 450804
rect 194501 450802 194567 450805
rect 191300 450800 194567 450802
rect 191300 450744 194506 450800
rect 194562 450744 194567 450800
rect 191300 450742 194567 450744
rect 191300 450740 191306 450742
rect 194501 450739 194567 450742
rect 372429 450802 372495 450805
rect 408309 450802 408375 450805
rect 372429 450800 408375 450802
rect 372429 450744 372434 450800
rect 372490 450744 408314 450800
rect 408370 450744 408375 450800
rect 372429 450742 408375 450744
rect 372429 450739 372495 450742
rect 408309 450739 408375 450742
rect 192334 450604 192340 450668
rect 192404 450666 192410 450668
rect 298921 450666 298987 450669
rect 192404 450664 298987 450666
rect 192404 450608 298926 450664
rect 298982 450608 298987 450664
rect 192404 450606 298987 450608
rect 192404 450604 192410 450606
rect 298921 450603 298987 450606
rect 372521 450666 372587 450669
rect 408125 450666 408191 450669
rect 372521 450664 408191 450666
rect 372521 450608 372526 450664
rect 372582 450608 408130 450664
rect 408186 450608 408191 450664
rect 372521 450606 408191 450608
rect 372521 450603 372587 450606
rect 408125 450603 408191 450606
rect 191414 450468 191420 450532
rect 191484 450530 191490 450532
rect 194317 450530 194383 450533
rect 191484 450528 194383 450530
rect 191484 450472 194322 450528
rect 194378 450472 194383 450528
rect 191484 450470 194383 450472
rect 191484 450468 191490 450470
rect 194317 450467 194383 450470
rect 194501 450530 194567 450533
rect 316585 450530 316651 450533
rect 194501 450528 316651 450530
rect 194501 450472 194506 450528
rect 194562 450472 316590 450528
rect 316646 450472 316651 450528
rect 194501 450470 316651 450472
rect 194501 450467 194567 450470
rect 316585 450467 316651 450470
rect 320633 450530 320699 450533
rect 388437 450530 388503 450533
rect 320633 450528 388503 450530
rect 320633 450472 320638 450528
rect 320694 450472 388442 450528
rect 388498 450472 388503 450528
rect 320633 450470 388503 450472
rect 320633 450467 320699 450470
rect 388437 450467 388503 450470
rect 187366 450332 187372 450396
rect 187436 450394 187442 450396
rect 329833 450394 329899 450397
rect 187436 450392 329899 450394
rect 187436 450336 329838 450392
rect 329894 450336 329899 450392
rect 187436 450334 329899 450336
rect 187436 450332 187442 450334
rect 329833 450331 329899 450334
rect 340505 450394 340571 450397
rect 405457 450394 405523 450397
rect 340505 450392 405523 450394
rect 340505 450336 340510 450392
rect 340566 450336 405462 450392
rect 405518 450336 405523 450392
rect 340505 450334 405523 450336
rect 340505 450331 340571 450334
rect 405457 450331 405523 450334
rect 193806 450196 193812 450260
rect 193876 450258 193882 450260
rect 194133 450258 194199 450261
rect 193876 450256 194199 450258
rect 193876 450200 194138 450256
rect 194194 450200 194199 450256
rect 193876 450198 194199 450200
rect 193876 450196 193882 450198
rect 194133 450195 194199 450198
rect 194317 450258 194383 450261
rect 357433 450258 357499 450261
rect 194317 450256 357499 450258
rect 194317 450200 194322 450256
rect 194378 450200 357438 450256
rect 357494 450200 357499 450256
rect 194317 450198 357499 450200
rect 194317 450195 194383 450198
rect 357433 450195 357499 450198
rect 184657 450122 184723 450125
rect 354489 450122 354555 450125
rect 184657 450120 354555 450122
rect 184657 450064 184662 450120
rect 184718 450064 354494 450120
rect 354550 450064 354555 450120
rect 184657 450062 354555 450064
rect 184657 450059 184723 450062
rect 354489 450059 354555 450062
rect 14549 449986 14615 449989
rect 233417 449986 233483 449989
rect 14549 449984 233483 449986
rect 14549 449928 14554 449984
rect 14610 449928 233422 449984
rect 233478 449928 233483 449984
rect 14549 449926 233483 449928
rect 14549 449923 14615 449926
rect 233417 449923 233483 449926
rect 304809 449986 304875 449989
rect 388713 449986 388779 449989
rect 304809 449984 388779 449986
rect 304809 449928 304814 449984
rect 304870 449928 388718 449984
rect 388774 449928 388779 449984
rect 304809 449926 388779 449928
rect 304809 449923 304875 449926
rect 388713 449923 388779 449926
rect 18597 449850 18663 449853
rect 230473 449850 230539 449853
rect 18597 449848 230539 449850
rect 18597 449792 18602 449848
rect 18658 449792 230478 449848
rect 230534 449792 230539 449848
rect 18597 449790 230539 449792
rect 18597 449787 18663 449790
rect 230473 449787 230539 449790
rect 367001 449850 367067 449853
rect 416078 449850 416084 449852
rect 367001 449848 416084 449850
rect 367001 449792 367006 449848
rect 367062 449792 416084 449848
rect 367001 449790 416084 449792
rect 367001 449787 367067 449790
rect 416078 449788 416084 449790
rect 416148 449788 416154 449852
rect -960 449578 480 449668
rect 190126 449652 190132 449716
rect 190196 449714 190202 449716
rect 261385 449714 261451 449717
rect 190196 449712 261451 449714
rect 190196 449656 261390 449712
rect 261446 449656 261451 449712
rect 190196 449654 261451 449656
rect 190196 449652 190202 449654
rect 261385 449651 261451 449654
rect 383929 449714 383995 449717
rect 389214 449714 389220 449716
rect 383929 449712 389220 449714
rect 383929 449656 383934 449712
rect 383990 449656 389220 449712
rect 383929 449654 389220 449656
rect 383929 449651 383995 449654
rect 389214 449652 389220 449654
rect 389284 449652 389290 449716
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 387609 449578 387675 449581
rect 387609 449576 393330 449578
rect 387609 449520 387614 449576
rect 387670 449520 393330 449576
rect 387609 449518 393330 449520
rect 387609 449515 387675 449518
rect 194041 449308 194107 449309
rect 193990 449306 193996 449308
rect 193950 449246 193996 449306
rect 194060 449304 194107 449308
rect 194102 449248 194107 449304
rect 193990 449244 193996 449246
rect 194060 449244 194107 449248
rect 194041 449243 194107 449244
rect 393270 449170 393330 449518
rect 417550 449170 417556 449172
rect 393270 449110 417556 449170
rect 417550 449108 417556 449110
rect 417620 449108 417626 449172
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580809 431626 580875 431629
rect 583520 431626 584960 431716
rect 580809 431624 584960 431626
rect 580809 431568 580814 431624
rect 580870 431568 584960 431624
rect 580809 431566 584960 431568
rect 580809 431563 580875 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect -960 423542 674 423602
rect -960 423466 480 423542
rect 614 423466 674 423542
rect -960 423452 674 423466
rect 246 423406 674 423452
rect 246 422922 306 423406
rect 246 422862 6930 422922
rect 6870 422378 6930 422862
rect 191833 422378 191899 422381
rect 6870 422376 191899 422378
rect 6870 422320 191838 422376
rect 191894 422320 191899 422376
rect 6870 422318 191899 422320
rect 191833 422315 191899 422318
rect 191465 419658 191531 419661
rect 191833 419658 191899 419661
rect 191465 419656 191899 419658
rect 191465 419600 191470 419656
rect 191526 419600 191838 419656
rect 191894 419600 191899 419656
rect 191465 419598 191899 419600
rect 191465 419595 191531 419598
rect 191833 419595 191899 419598
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3693 410546 3759 410549
rect -960 410544 3759 410546
rect -960 410488 3698 410544
rect 3754 410488 3759 410544
rect -960 410486 3759 410488
rect -960 410396 480 410486
rect 3693 410483 3759 410486
rect 580901 404970 580967 404973
rect 583520 404970 584960 405060
rect 580901 404968 584960 404970
rect 580901 404912 580906 404968
rect 580962 404912 584960 404968
rect 580901 404910 584960 404912
rect 580901 404907 580967 404910
rect 583520 404820 584960 404910
rect 190821 398850 190887 398853
rect 191097 398850 191163 398853
rect 190821 398848 191163 398850
rect 190821 398792 190826 398848
rect 190882 398792 191102 398848
rect 191158 398792 191163 398848
rect 190821 398790 191163 398792
rect 190821 398787 190887 398790
rect 191097 398787 191163 398790
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 190821 397354 190887 397357
rect 191097 397354 191163 397357
rect 190821 397352 191163 397354
rect 190821 397296 190826 397352
rect 190882 397296 191102 397352
rect 191158 397296 191163 397352
rect 190821 397294 191163 397296
rect 190821 397291 190887 397294
rect 191097 397291 191163 397294
rect 191465 397354 191531 397357
rect 191833 397354 191899 397357
rect 191465 397352 191899 397354
rect 191465 397296 191470 397352
rect 191526 397296 191838 397352
rect 191894 397296 191899 397352
rect 191465 397294 191899 397296
rect 191465 397291 191531 397294
rect 191833 397291 191899 397294
rect 191833 395994 191899 395997
rect 192334 395994 192340 395996
rect 191833 395992 192340 395994
rect 191833 395936 191838 395992
rect 191894 395936 192340 395992
rect 191833 395934 192340 395936
rect 191833 395931 191899 395934
rect 192334 395932 192340 395934
rect 192404 395932 192410 395996
rect 186773 394770 186839 394773
rect 192334 394770 192340 394772
rect 186773 394768 192340 394770
rect 186773 394712 186778 394768
rect 186834 394712 192340 394768
rect 186773 394710 192340 394712
rect 186773 394707 186839 394710
rect 192334 394708 192340 394710
rect 192404 394708 192410 394772
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 190821 372602 190887 372605
rect 191373 372602 191439 372605
rect 190821 372600 191439 372602
rect 190821 372544 190826 372600
rect 190882 372544 191378 372600
rect 191434 372544 191439 372600
rect 190821 372542 191439 372544
rect 190821 372539 190887 372542
rect 191373 372539 191439 372542
rect -960 371378 480 371468
rect 3049 371378 3115 371381
rect -960 371376 3115 371378
rect -960 371320 3054 371376
rect 3110 371320 3115 371376
rect -960 371318 3115 371320
rect -960 371228 480 371318
rect 3049 371315 3115 371318
rect 191373 369882 191439 369885
rect 192150 369882 192156 369884
rect 191373 369880 192156 369882
rect 191373 369824 191378 369880
rect 191434 369824 192156 369880
rect 191373 369822 192156 369824
rect 191373 369819 191439 369822
rect 192150 369820 192156 369822
rect 192220 369820 192226 369884
rect 191833 369204 191899 369205
rect 191782 369202 191788 369204
rect 191742 369142 191788 369202
rect 191852 369200 191899 369204
rect 191894 369144 191899 369200
rect 191782 369140 191788 369142
rect 191852 369140 191899 369144
rect 191833 369139 191899 369140
rect 188153 369066 188219 369069
rect 191833 369066 191899 369069
rect 188153 369064 191899 369066
rect 188153 369008 188158 369064
rect 188214 369008 191838 369064
rect 191894 369008 191899 369064
rect 188153 369006 191899 369008
rect 188153 369003 188219 369006
rect 191833 369003 191899 369006
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2957 319290 3023 319293
rect -960 319288 3023 319290
rect -960 319232 2962 319288
rect 3018 319232 3023 319288
rect -960 319230 3023 319232
rect -960 319140 480 319230
rect 2957 319227 3023 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580809 298754 580875 298757
rect 583520 298754 584960 298844
rect 580809 298752 584960 298754
rect 580809 298696 580814 298752
rect 580870 298696 584960 298752
rect 580809 298694 584960 298696
rect 580809 298691 580875 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 2865 293178 2931 293181
rect -960 293176 2931 293178
rect -960 293120 2870 293176
rect 2926 293120 2931 293176
rect -960 293118 2931 293120
rect -960 293028 480 293118
rect 2865 293115 2931 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 190126 249052 190132 249116
rect 190196 249114 190202 249116
rect 217317 249114 217383 249117
rect 190196 249112 217383 249114
rect 190196 249056 217322 249112
rect 217378 249056 217383 249112
rect 190196 249054 217383 249056
rect 190196 249052 190202 249054
rect 217317 249051 217383 249054
rect 201677 248298 201743 248301
rect 226425 248298 226491 248301
rect 201677 248296 226491 248298
rect 201677 248240 201682 248296
rect 201738 248240 226430 248296
rect 226486 248240 226491 248296
rect 201677 248238 226491 248240
rect 201677 248235 201743 248238
rect 226425 248235 226491 248238
rect 222837 248162 222903 248165
rect 254025 248162 254091 248165
rect 222837 248160 254091 248162
rect 222837 248104 222842 248160
rect 222898 248104 254030 248160
rect 254086 248104 254091 248160
rect 222837 248102 254091 248104
rect 222837 248099 222903 248102
rect 254025 248099 254091 248102
rect 214557 248026 214623 248029
rect 223665 248026 223731 248029
rect 214557 248024 223731 248026
rect 214557 247968 214562 248024
rect 214618 247968 223670 248024
rect 223726 247968 223731 248024
rect 214557 247966 223731 247968
rect 214557 247963 214623 247966
rect 223665 247963 223731 247966
rect 225781 248026 225847 248029
rect 258165 248026 258231 248029
rect 225781 248024 258231 248026
rect 225781 247968 225786 248024
rect 225842 247968 258170 248024
rect 258226 247968 258231 248024
rect 225781 247966 258231 247968
rect 225781 247963 225847 247966
rect 258165 247963 258231 247966
rect 347865 248026 347931 248029
rect 358077 248026 358143 248029
rect 347865 248024 358143 248026
rect 347865 247968 347870 248024
rect 347926 247968 358082 248024
rect 358138 247968 358143 248024
rect 347865 247966 358143 247968
rect 347865 247963 347931 247966
rect 358077 247963 358143 247966
rect 213177 247890 213243 247893
rect 222285 247890 222351 247893
rect 213177 247888 222351 247890
rect 213177 247832 213182 247888
rect 213238 247832 222290 247888
rect 222346 247832 222351 247888
rect 213177 247830 222351 247832
rect 213177 247827 213243 247830
rect 222285 247827 222351 247830
rect 223021 247890 223087 247893
rect 256785 247890 256851 247893
rect 223021 247888 256851 247890
rect 223021 247832 223026 247888
rect 223082 247832 256790 247888
rect 256846 247832 256851 247888
rect 223021 247830 256851 247832
rect 223021 247827 223087 247830
rect 256785 247827 256851 247830
rect 343725 247890 343791 247893
rect 356789 247890 356855 247893
rect 343725 247888 356855 247890
rect 343725 247832 343730 247888
rect 343786 247832 356794 247888
rect 356850 247832 356855 247888
rect 343725 247830 356855 247832
rect 343725 247827 343791 247830
rect 356789 247827 356855 247830
rect 197353 247754 197419 247757
rect 225045 247754 225111 247757
rect 197353 247752 225111 247754
rect 197353 247696 197358 247752
rect 197414 247696 225050 247752
rect 225106 247696 225111 247752
rect 197353 247694 225111 247696
rect 197353 247691 197419 247694
rect 225045 247691 225111 247694
rect 225597 247754 225663 247757
rect 260925 247754 260991 247757
rect 225597 247752 260991 247754
rect 225597 247696 225602 247752
rect 225658 247696 260930 247752
rect 260986 247696 260991 247752
rect 225597 247694 260991 247696
rect 225597 247691 225663 247694
rect 260925 247691 260991 247694
rect 345105 247754 345171 247757
rect 358261 247754 358327 247757
rect 345105 247752 358327 247754
rect 345105 247696 345110 247752
rect 345166 247696 358266 247752
rect 358322 247696 358327 247752
rect 345105 247694 358327 247696
rect 345105 247691 345171 247694
rect 358261 247691 358327 247694
rect 186313 247618 186379 247621
rect 220905 247618 220971 247621
rect 186313 247616 220971 247618
rect 186313 247560 186318 247616
rect 186374 247560 220910 247616
rect 220966 247560 220971 247616
rect 186313 247558 220971 247560
rect 186313 247555 186379 247558
rect 220905 247555 220971 247558
rect 228357 247618 228423 247621
rect 265065 247618 265131 247621
rect 228357 247616 265131 247618
rect 228357 247560 228362 247616
rect 228418 247560 265070 247616
rect 265126 247560 265131 247616
rect 228357 247558 265131 247560
rect 228357 247555 228423 247558
rect 265065 247555 265131 247558
rect 340965 247618 341031 247621
rect 360837 247618 360903 247621
rect 340965 247616 360903 247618
rect 340965 247560 340970 247616
rect 341026 247560 360842 247616
rect 360898 247560 360903 247616
rect 340965 247558 360903 247560
rect 340965 247555 341031 247558
rect 360837 247555 360903 247558
rect 208393 247482 208459 247485
rect 229185 247482 229251 247485
rect 208393 247480 229251 247482
rect 208393 247424 208398 247480
rect 208454 247424 229190 247480
rect 229246 247424 229251 247480
rect 208393 247422 229251 247424
rect 208393 247419 208459 247422
rect 229185 247419 229251 247422
rect 215937 247346 216003 247349
rect 227805 247346 227871 247349
rect 215937 247344 227871 247346
rect 215937 247288 215942 247344
rect 215998 247288 227810 247344
rect 227866 247288 227871 247344
rect 215937 247286 227871 247288
rect 215937 247283 216003 247286
rect 227805 247283 227871 247286
rect 353385 247346 353451 247349
rect 357157 247346 357223 247349
rect 353385 247344 357223 247346
rect 353385 247288 353390 247344
rect 353446 247288 357162 247344
rect 357218 247288 357223 247344
rect 353385 247286 357223 247288
rect 353385 247283 353451 247286
rect 357157 247283 357223 247286
rect 356145 247210 356211 247213
rect 357198 247210 357204 247212
rect 356145 247208 357204 247210
rect 356145 247152 356150 247208
rect 356206 247152 357204 247208
rect 356145 247150 357204 247152
rect 356145 247147 356211 247150
rect 357198 247148 357204 247150
rect 357268 247148 357274 247212
rect 354765 247074 354831 247077
rect 356973 247074 357039 247077
rect 354765 247072 357039 247074
rect 354765 247016 354770 247072
rect 354826 247016 356978 247072
rect 357034 247016 357039 247072
rect 354765 247014 357039 247016
rect 354765 247011 354831 247014
rect 356973 247011 357039 247014
rect 358905 247074 358971 247077
rect 359958 247074 359964 247076
rect 358905 247072 359964 247074
rect 358905 247016 358910 247072
rect 358966 247016 359964 247072
rect 358905 247014 359964 247016
rect 358905 247011 358971 247014
rect 359958 247012 359964 247014
rect 360028 247012 360034 247076
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 580717 232386 580783 232389
rect 583520 232386 584960 232476
rect 580717 232384 584960 232386
rect 580717 232328 580722 232384
rect 580778 232328 584960 232384
rect 580717 232326 584960 232328
rect 580717 232323 580783 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580625 219058 580691 219061
rect 583520 219058 584960 219148
rect 580625 219056 584960 219058
rect 580625 219000 580630 219056
rect 580686 219000 584960 219056
rect 580625 218998 584960 219000
rect 580625 218995 580691 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 150985 196076 151051 196077
rect 551001 196076 551067 196077
rect 150934 196074 150940 196076
rect 150894 196014 150940 196074
rect 151004 196072 151051 196076
rect 550950 196074 550956 196076
rect 151046 196016 151051 196072
rect 150934 196012 150940 196014
rect 151004 196012 151051 196016
rect 550910 196014 550956 196074
rect 551020 196072 551067 196076
rect 551062 196016 551067 196072
rect 550950 196012 550956 196014
rect 551020 196012 551067 196016
rect 150985 196011 151051 196012
rect 551001 196011 551067 196012
rect 193990 193972 193996 194036
rect 194060 194034 194066 194036
rect 580809 194034 580875 194037
rect 194060 194032 580875 194034
rect 194060 193976 580814 194032
rect 580870 193976 580875 194032
rect 194060 193974 580875 193976
rect 194060 193972 194066 193974
rect 580809 193971 580875 193974
rect 193806 193836 193812 193900
rect 193876 193898 193882 193900
rect 580625 193898 580691 193901
rect 193876 193896 580691 193898
rect 193876 193840 580630 193896
rect 580686 193840 580691 193896
rect 193876 193838 580691 193840
rect 193876 193836 193882 193838
rect 580625 193835 580691 193838
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect 158713 189274 158779 189277
rect 156558 189272 158779 189274
rect 156558 189216 158718 189272
rect 158774 189216 158779 189272
rect 156558 189214 158779 189216
rect 156558 189190 156618 189214
rect 158713 189211 158779 189214
rect 556570 189138 556630 189190
rect 558913 189138 558979 189141
rect 556570 189136 558979 189138
rect 556570 189080 558918 189136
rect 558974 189080 558979 189136
rect 556570 189078 558979 189080
rect 558913 189075 558979 189078
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 580441 179210 580507 179213
rect 583520 179210 584960 179300
rect 580441 179208 584960 179210
rect 580441 179152 580446 179208
rect 580502 179152 584960 179208
rect 580441 179150 584960 179152
rect 580441 179147 580507 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3601 162890 3667 162893
rect -960 162888 3667 162890
rect -960 162832 3606 162888
rect 3662 162832 3667 162888
rect -960 162830 3667 162832
rect -960 162740 480 162830
rect 3601 162827 3667 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3785 149834 3851 149837
rect -960 149832 3851 149834
rect -960 149776 3790 149832
rect 3846 149776 3851 149832
rect -960 149774 3851 149776
rect -960 149684 480 149774
rect 3785 149771 3851 149774
rect 16757 146978 16823 146981
rect 17309 146978 17375 146981
rect 416773 146978 416839 146981
rect 417325 146978 417391 146981
rect 16757 146976 19442 146978
rect 16757 146920 16762 146976
rect 16818 146920 17314 146976
rect 17370 146924 19442 146976
rect 416773 146976 419458 146978
rect 17370 146920 20056 146924
rect 16757 146918 20056 146920
rect 16757 146915 16823 146918
rect 17309 146915 17375 146918
rect 19382 146864 20056 146918
rect 416773 146920 416778 146976
rect 416834 146920 417330 146976
rect 417386 146924 419458 146976
rect 417386 146920 420072 146924
rect 416773 146918 420072 146920
rect 416773 146915 416839 146918
rect 417325 146915 417391 146918
rect 419398 146864 420072 146918
rect 17401 146026 17467 146029
rect 17677 146026 17743 146029
rect 17401 146024 19442 146026
rect 17401 145968 17406 146024
rect 17462 145968 17682 146024
rect 17738 145972 19442 146024
rect 17738 145968 20056 145972
rect 17401 145966 20056 145968
rect 17401 145963 17467 145966
rect 17677 145963 17743 145966
rect 19382 145912 20056 145966
rect 417182 145964 417188 146028
rect 417252 146026 417258 146028
rect 417734 146026 417740 146028
rect 417252 145966 417740 146026
rect 417252 145964 417258 145966
rect 417734 145964 417740 145966
rect 417804 146026 417810 146028
rect 417804 145972 419458 146026
rect 417804 145966 420072 145972
rect 417804 145964 417810 145966
rect 419398 145912 420072 145966
rect 16941 144802 17007 144805
rect 17677 144802 17743 144805
rect 16941 144800 17743 144802
rect 16941 144744 16946 144800
rect 17002 144744 17682 144800
rect 17738 144744 17743 144800
rect 16941 144742 17743 144744
rect 16941 144739 17007 144742
rect 17677 144739 17743 144742
rect 17677 143850 17743 143853
rect 417141 143850 417207 143853
rect 17677 143848 19442 143850
rect 17677 143792 17682 143848
rect 17738 143796 19442 143848
rect 417141 143848 419458 143850
rect 17738 143792 20056 143796
rect 17677 143790 20056 143792
rect 17677 143787 17743 143790
rect 19382 143736 20056 143790
rect 417141 143792 417146 143848
rect 417202 143796 419458 143848
rect 417202 143792 420072 143796
rect 417141 143790 420072 143792
rect 417141 143787 417207 143790
rect 419398 143736 420072 143790
rect 17585 142898 17651 142901
rect 17585 142896 19442 142898
rect 17585 142840 17590 142896
rect 17646 142844 19442 142896
rect 17646 142840 20056 142844
rect 17585 142838 20056 142840
rect 17585 142835 17651 142838
rect 19382 142784 20056 142838
rect 419398 142784 420072 142844
rect 390185 142762 390251 142765
rect 417734 142762 417740 142764
rect 390185 142760 417740 142762
rect 390185 142704 390190 142760
rect 390246 142704 417740 142760
rect 390185 142702 417740 142704
rect 390185 142699 390251 142702
rect 417734 142700 417740 142702
rect 417804 142762 417810 142764
rect 419398 142762 419458 142784
rect 417804 142702 419458 142762
rect 417804 142700 417810 142702
rect 416773 141130 416839 141133
rect 417509 141130 417575 141133
rect 416773 141128 419458 141130
rect 19382 141016 20056 141076
rect 416773 141072 416778 141128
rect 416834 141072 417514 141128
rect 417570 141076 419458 141128
rect 417570 141072 420072 141076
rect 416773 141070 420072 141072
rect 416773 141067 416839 141070
rect 417509 141067 417575 141070
rect 419398 141016 420072 141070
rect 16849 140858 16915 140861
rect 17769 140858 17835 140861
rect 19382 140858 19442 141016
rect 16849 140856 19442 140858
rect 16849 140800 16854 140856
rect 16910 140800 17774 140856
rect 17830 140800 19442 140856
rect 16849 140798 19442 140800
rect 16849 140795 16915 140798
rect 17769 140795 17835 140798
rect 16665 140042 16731 140045
rect 17585 140042 17651 140045
rect 416773 140042 416839 140045
rect 417233 140042 417299 140045
rect 16665 140040 19442 140042
rect 16665 139984 16670 140040
rect 16726 139984 17590 140040
rect 17646 139988 19442 140040
rect 416773 140040 419458 140042
rect 17646 139984 20056 139988
rect 16665 139982 20056 139984
rect 16665 139979 16731 139982
rect 17585 139979 17651 139982
rect 19382 139928 20056 139982
rect 416773 139984 416778 140040
rect 416834 139984 417238 140040
rect 417294 139988 419458 140040
rect 417294 139984 420072 139988
rect 416773 139982 420072 139984
rect 416773 139979 416839 139982
rect 417233 139979 417299 139982
rect 419398 139928 420072 139982
rect 580533 139362 580599 139365
rect 583520 139362 584960 139452
rect 580533 139360 584960 139362
rect 580533 139304 580538 139360
rect 580594 139304 584960 139360
rect 580533 139302 584960 139304
rect 580533 139299 580599 139302
rect 583520 139212 584960 139302
rect 17861 138274 17927 138277
rect 17861 138272 19442 138274
rect 17861 138216 17866 138272
rect 17922 138220 19442 138272
rect 17922 138216 20056 138220
rect 17861 138214 20056 138216
rect 17861 138211 17927 138214
rect 19382 138160 20056 138214
rect 417550 138212 417556 138276
rect 417620 138274 417626 138276
rect 417918 138274 417924 138276
rect 417620 138214 417924 138274
rect 417620 138212 417626 138214
rect 417918 138212 417924 138214
rect 417988 138274 417994 138276
rect 417988 138220 419458 138274
rect 417988 138214 420072 138220
rect 417988 138212 417994 138214
rect 419398 138160 420072 138214
rect -960 136778 480 136868
rect 3049 136778 3115 136781
rect -960 136776 3115 136778
rect -960 136720 3054 136776
rect 3110 136720 3115 136776
rect -960 136718 3115 136720
rect -960 136628 480 136718
rect 3049 136715 3115 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 17033 120050 17099 120053
rect 417141 120050 417207 120053
rect 17033 120048 19442 120050
rect 17033 119992 17038 120048
rect 17094 119996 19442 120048
rect 417141 120048 419458 120050
rect 17094 119992 20056 119996
rect 17033 119990 20056 119992
rect 17033 119987 17099 119990
rect 19382 119936 20056 119990
rect 417141 119992 417146 120048
rect 417202 119996 419458 120048
rect 417202 119992 420072 119996
rect 417141 119990 420072 119992
rect 417141 119987 417207 119990
rect 419398 119936 420072 119990
rect 17217 118418 17283 118421
rect 417785 118418 417851 118421
rect 17217 118416 19442 118418
rect 17217 118360 17222 118416
rect 17278 118364 19442 118416
rect 417785 118416 419458 118418
rect 17278 118360 20056 118364
rect 17217 118358 20056 118360
rect 17217 118355 17283 118358
rect 19382 118304 20056 118358
rect 417785 118360 417790 118416
rect 417846 118364 419458 118416
rect 417846 118360 420072 118364
rect 417785 118358 420072 118360
rect 417785 118355 417851 118358
rect 419398 118304 420072 118358
rect 18781 118146 18847 118149
rect 417417 118146 417483 118149
rect 18781 118144 19442 118146
rect 18781 118088 18786 118144
rect 18842 118092 19442 118144
rect 417417 118144 419458 118146
rect 18842 118088 20056 118092
rect 18781 118086 20056 118088
rect 18781 118083 18847 118086
rect 19382 118032 20056 118086
rect 417417 118088 417422 118144
rect 417478 118092 419458 118144
rect 417478 118088 420072 118092
rect 417417 118086 420072 118088
rect 417417 118083 417483 118086
rect 419398 118032 420072 118086
rect 579981 112842 580047 112845
rect 583520 112842 584960 112932
rect 579981 112840 584960 112842
rect 579981 112784 579986 112840
rect 580042 112784 584960 112840
rect 579981 112782 584960 112784
rect 579981 112779 580047 112782
rect 583520 112692 584960 112782
rect 342253 111210 342319 111213
rect 419758 111210 419764 111212
rect 342253 111208 419764 111210
rect 342253 111152 342258 111208
rect 342314 111152 419764 111208
rect 342253 111150 419764 111152
rect 342253 111147 342319 111150
rect 419758 111148 419764 111150
rect 419828 111148 419834 111212
rect 336733 111074 336799 111077
rect 419942 111074 419948 111076
rect 336733 111072 419948 111074
rect 336733 111016 336738 111072
rect 336794 111016 419948 111072
rect 336733 111014 419948 111016
rect 336733 111011 336799 111014
rect 419942 111012 419948 111014
rect 420012 111012 420018 111076
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 451273 109852 451339 109853
rect 480897 109852 480963 109853
rect 483473 109852 483539 109853
rect 485957 109852 486023 109853
rect 488257 109852 488323 109853
rect 491017 109852 491083 109853
rect 451273 109848 451286 109852
rect 451350 109850 451356 109852
rect 451273 109792 451278 109848
rect 451273 109788 451286 109792
rect 451350 109790 451430 109850
rect 480897 109848 480934 109852
rect 480998 109850 481004 109852
rect 480897 109792 480902 109848
rect 451350 109788 451356 109790
rect 480897 109788 480934 109792
rect 480998 109790 481054 109850
rect 483473 109848 483518 109852
rect 483582 109850 483588 109852
rect 483473 109792 483478 109848
rect 480998 109788 481004 109790
rect 483473 109788 483518 109792
rect 483582 109790 483630 109850
rect 485957 109848 485966 109852
rect 486030 109850 486036 109852
rect 485957 109792 485962 109848
rect 483582 109788 483588 109790
rect 485957 109788 485966 109792
rect 486030 109790 486114 109850
rect 488257 109848 488278 109852
rect 488342 109850 488348 109852
rect 490992 109850 490998 109852
rect 488257 109792 488262 109848
rect 486030 109788 486036 109790
rect 488257 109788 488278 109792
rect 488342 109790 488414 109850
rect 490926 109790 490998 109850
rect 491062 109848 491083 109852
rect 491078 109792 491083 109848
rect 488342 109788 488348 109790
rect 490992 109788 490998 109790
rect 491062 109788 491083 109792
rect 451273 109787 451339 109788
rect 480897 109787 480963 109788
rect 483473 109787 483539 109788
rect 485957 109787 486023 109788
rect 488257 109787 488323 109788
rect 491017 109787 491083 109788
rect 476113 109716 476179 109717
rect 476062 109714 476068 109716
rect 476022 109654 476068 109714
rect 476132 109712 476179 109716
rect 476174 109656 476179 109712
rect 476062 109652 476068 109654
rect 476132 109652 476179 109656
rect 476113 109651 476179 109652
rect 493409 109716 493475 109717
rect 495893 109716 495959 109717
rect 498469 109716 498535 109717
rect 493409 109712 493446 109716
rect 493510 109714 493516 109716
rect 495888 109714 495894 109716
rect 493409 109656 493414 109712
rect 493409 109652 493446 109656
rect 493510 109654 493566 109714
rect 495802 109654 495894 109714
rect 493510 109652 493516 109654
rect 495888 109652 495894 109654
rect 495958 109652 495964 109716
rect 498469 109712 498478 109716
rect 498542 109714 498548 109716
rect 498469 109656 498474 109712
rect 498469 109652 498478 109656
rect 498542 109654 498626 109714
rect 498542 109652 498548 109654
rect 493409 109651 493475 109652
rect 495893 109651 495959 109652
rect 498469 109651 498535 109652
rect 50797 109580 50863 109581
rect 56041 109580 56107 109581
rect 61101 109580 61167 109581
rect 105997 109580 106063 109581
rect 108573 109580 108639 109581
rect 50736 109578 50742 109580
rect 50706 109518 50742 109578
rect 50806 109576 50863 109580
rect 50858 109520 50863 109576
rect 50736 109516 50742 109518
rect 50806 109516 50863 109520
rect 56040 109516 56046 109580
rect 56110 109578 56116 109580
rect 61072 109578 61078 109580
rect 56110 109518 56198 109578
rect 61010 109518 61078 109578
rect 61142 109576 61167 109580
rect 105952 109578 105958 109580
rect 61162 109520 61167 109576
rect 56110 109516 56116 109518
rect 61072 109516 61078 109518
rect 61142 109516 61167 109520
rect 105906 109518 105958 109578
rect 106022 109576 106063 109580
rect 108536 109578 108542 109580
rect 106058 109520 106063 109576
rect 105952 109516 105958 109518
rect 106022 109516 106063 109520
rect 108482 109518 108542 109578
rect 108606 109576 108639 109580
rect 108634 109520 108639 109576
rect 108536 109516 108542 109518
rect 108606 109516 108639 109520
rect 50797 109515 50863 109516
rect 56041 109515 56107 109516
rect 61101 109515 61167 109516
rect 105997 109515 106063 109516
rect 108573 109515 108639 109516
rect 456977 109580 457043 109581
rect 505921 109580 505987 109581
rect 508497 109580 508563 109581
rect 515857 109580 515923 109581
rect 518433 109580 518499 109581
rect 456977 109576 456998 109580
rect 457062 109578 457068 109580
rect 456977 109520 456982 109576
rect 456977 109516 456998 109520
rect 457062 109518 457134 109578
rect 457062 109516 457068 109518
rect 461072 109516 461078 109580
rect 461142 109516 461148 109580
rect 505921 109576 505958 109580
rect 506022 109578 506028 109580
rect 505921 109520 505926 109576
rect 505921 109516 505958 109520
rect 506022 109518 506078 109578
rect 508497 109576 508542 109580
rect 508606 109578 508612 109580
rect 508497 109520 508502 109576
rect 506022 109516 506028 109518
rect 508497 109516 508542 109520
rect 508606 109518 508654 109578
rect 515857 109576 515886 109580
rect 515950 109578 515956 109580
rect 515857 109520 515862 109576
rect 508606 109516 508612 109518
rect 515857 109516 515886 109520
rect 515950 109518 516014 109578
rect 518433 109576 518470 109580
rect 518534 109578 518540 109580
rect 518433 109520 518438 109576
rect 515950 109516 515956 109518
rect 518433 109516 518470 109520
rect 518534 109518 518590 109578
rect 518534 109516 518540 109518
rect 456977 109515 457043 109516
rect 408309 109306 408375 109309
rect 461080 109306 461140 109516
rect 505921 109515 505987 109516
rect 508497 109515 508563 109516
rect 515857 109515 515923 109516
rect 518433 109515 518499 109516
rect 408309 109304 461140 109306
rect 408309 109248 408314 109304
rect 408370 109248 461140 109304
rect 408309 109246 461140 109248
rect 408309 109243 408375 109246
rect 407665 109170 407731 109173
rect 468334 109170 468340 109172
rect 407665 109168 468340 109170
rect 407665 109112 407670 109168
rect 407726 109112 468340 109168
rect 407665 109110 468340 109112
rect 407665 109107 407731 109110
rect 468334 109108 468340 109110
rect 468404 109108 468410 109172
rect 48313 109036 48379 109037
rect 68369 109036 68435 109037
rect 100937 109036 101003 109037
rect 111057 109036 111123 109037
rect 113449 109036 113515 109037
rect 48262 109034 48268 109036
rect 48222 108974 48268 109034
rect 48332 109032 48379 109036
rect 68318 109034 68324 109036
rect 48374 108976 48379 109032
rect 48262 108972 48268 108974
rect 48332 108972 48379 108976
rect 68278 108974 68324 109034
rect 68388 109032 68435 109036
rect 100886 109034 100892 109036
rect 68430 108976 68435 109032
rect 68318 108972 68324 108974
rect 68388 108972 68435 108976
rect 100846 108974 100892 109034
rect 100956 109032 101003 109036
rect 111006 109034 111012 109036
rect 100998 108976 101003 109032
rect 100886 108972 100892 108974
rect 100956 108972 101003 108976
rect 110966 108974 111012 109034
rect 111076 109032 111123 109036
rect 113398 109034 113404 109036
rect 111118 108976 111123 109032
rect 111006 108972 111012 108974
rect 111076 108972 111123 108976
rect 113358 108974 113404 109034
rect 113468 109032 113515 109036
rect 113510 108976 113515 109032
rect 113398 108972 113404 108974
rect 113468 108972 113515 108976
rect 125910 108972 125916 109036
rect 125980 109034 125986 109036
rect 389214 109034 389220 109036
rect 125980 108974 389220 109034
rect 125980 108972 125986 108974
rect 389214 108972 389220 108974
rect 389284 108972 389290 109036
rect 407849 109034 407915 109037
rect 500953 109036 501019 109037
rect 470910 109034 470916 109036
rect 407849 109032 470916 109034
rect 407849 108976 407854 109032
rect 407910 108976 470916 109032
rect 407849 108974 470916 108976
rect 48313 108971 48379 108972
rect 68369 108971 68435 108972
rect 100937 108971 101003 108972
rect 111057 108971 111123 108972
rect 113449 108971 113515 108972
rect 407849 108971 407915 108974
rect 470910 108972 470916 108974
rect 470980 108972 470986 109036
rect 500902 109034 500908 109036
rect 500862 108974 500908 109034
rect 500972 109032 501019 109036
rect 501014 108976 501019 109032
rect 500902 108972 500908 108974
rect 500972 108972 501019 108976
rect 500953 108971 501019 108972
rect 503437 109036 503503 109037
rect 513373 109036 513439 109037
rect 520917 109036 520983 109037
rect 523309 109036 523375 109037
rect 525885 109036 525951 109037
rect 503437 109032 503484 109036
rect 503548 109034 503554 109036
rect 503437 108976 503442 109032
rect 503437 108972 503484 108976
rect 503548 108974 503594 109034
rect 513373 109032 513420 109036
rect 513484 109034 513490 109036
rect 513373 108976 513378 109032
rect 503548 108972 503554 108974
rect 513373 108972 513420 108976
rect 513484 108974 513530 109034
rect 520917 109032 520964 109036
rect 521028 109034 521034 109036
rect 520917 108976 520922 109032
rect 513484 108972 513490 108974
rect 520917 108972 520964 108976
rect 521028 108974 521074 109034
rect 523309 109032 523356 109036
rect 523420 109034 523426 109036
rect 523309 108976 523314 109032
rect 521028 108972 521034 108974
rect 523309 108972 523356 108976
rect 523420 108974 523466 109034
rect 525885 109032 525932 109036
rect 525996 109034 526002 109036
rect 525885 108976 525890 109032
rect 523420 108972 523426 108974
rect 525885 108972 525932 108976
rect 525996 108974 526042 109034
rect 525996 108972 526002 108974
rect 503437 108971 503503 108972
rect 513373 108971 513439 108972
rect 520917 108971 520983 108972
rect 523309 108971 523375 108972
rect 525885 108971 525951 108972
rect 65926 108836 65932 108900
rect 65996 108898 66002 108900
rect 188470 108898 188476 108900
rect 65996 108838 188476 108898
rect 65996 108836 66002 108838
rect 188470 108836 188476 108838
rect 188540 108836 188546 108900
rect 408217 108898 408283 108901
rect 465942 108898 465948 108900
rect 408217 108896 465948 108898
rect 408217 108840 408222 108896
rect 408278 108840 465948 108896
rect 408217 108838 465948 108840
rect 408217 108835 408283 108838
rect 465942 108836 465948 108838
rect 466012 108836 466018 108900
rect 53649 108764 53715 108765
rect 53598 108762 53604 108764
rect 53558 108702 53604 108762
rect 53668 108760 53715 108764
rect 53710 108704 53715 108760
rect 53598 108700 53604 108702
rect 53668 108700 53715 108704
rect 90950 108700 90956 108764
rect 91020 108762 91026 108764
rect 186814 108762 186820 108764
rect 91020 108702 186820 108762
rect 91020 108700 91026 108702
rect 186814 108700 186820 108702
rect 186884 108700 186890 108764
rect 53649 108699 53715 108700
rect 95918 108564 95924 108628
rect 95988 108626 95994 108628
rect 187182 108626 187188 108628
rect 95988 108566 187188 108626
rect 95988 108564 95994 108566
rect 187182 108564 187188 108566
rect 187252 108564 187258 108628
rect 457989 108492 458055 108493
rect 118550 108428 118556 108492
rect 118620 108490 118626 108492
rect 184238 108490 184244 108492
rect 118620 108430 184244 108490
rect 118620 108428 118626 108430
rect 184238 108428 184244 108430
rect 184308 108428 184314 108492
rect 457989 108488 458036 108492
rect 458100 108490 458106 108492
rect 457989 108432 457994 108488
rect 457989 108428 458036 108432
rect 458100 108430 458146 108490
rect 458100 108428 458106 108430
rect 457989 108427 458055 108428
rect 19793 107538 19859 107541
rect 35893 107540 35959 107541
rect 19926 107538 19932 107540
rect 19793 107536 19932 107538
rect 19793 107480 19798 107536
rect 19854 107480 19932 107536
rect 19793 107478 19932 107480
rect 19793 107475 19859 107478
rect 19926 107476 19932 107478
rect 19996 107476 20002 107540
rect 35893 107536 35940 107540
rect 36004 107538 36010 107540
rect 36905 107538 36971 107541
rect 38101 107540 38167 107541
rect 39573 107540 39639 107541
rect 40493 107540 40559 107541
rect 43161 107540 43227 107541
rect 44265 107540 44331 107541
rect 45369 107540 45435 107541
rect 37038 107538 37044 107540
rect 35893 107480 35898 107536
rect 35893 107476 35940 107480
rect 36004 107478 36050 107538
rect 36905 107536 37044 107538
rect 36905 107480 36910 107536
rect 36966 107480 37044 107536
rect 36905 107478 37044 107480
rect 36004 107476 36010 107478
rect 35893 107475 35959 107476
rect 36905 107475 36971 107478
rect 37038 107476 37044 107478
rect 37108 107476 37114 107540
rect 38101 107536 38148 107540
rect 38212 107538 38218 107540
rect 38101 107480 38106 107536
rect 38101 107476 38148 107480
rect 38212 107478 38258 107538
rect 39573 107536 39620 107540
rect 39684 107538 39690 107540
rect 39573 107480 39578 107536
rect 38212 107476 38218 107478
rect 39573 107476 39620 107480
rect 39684 107478 39730 107538
rect 40493 107536 40540 107540
rect 40604 107538 40610 107540
rect 43110 107538 43116 107540
rect 40493 107480 40498 107536
rect 39684 107476 39690 107478
rect 40493 107476 40540 107480
rect 40604 107478 40650 107538
rect 43070 107478 43116 107538
rect 43180 107536 43227 107540
rect 44214 107538 44220 107540
rect 43222 107480 43227 107536
rect 40604 107476 40610 107478
rect 43110 107476 43116 107478
rect 43180 107476 43227 107480
rect 44174 107478 44220 107538
rect 44284 107536 44331 107540
rect 45318 107538 45324 107540
rect 44326 107480 44331 107536
rect 44214 107476 44220 107478
rect 44284 107476 44331 107480
rect 45278 107478 45324 107538
rect 45388 107536 45435 107540
rect 45430 107480 45435 107536
rect 45318 107476 45324 107478
rect 45388 107476 45435 107480
rect 38101 107475 38167 107476
rect 39573 107475 39639 107476
rect 40493 107475 40559 107476
rect 43161 107475 43227 107476
rect 44265 107475 44331 107476
rect 45369 107475 45435 107476
rect 46565 107540 46631 107541
rect 47577 107540 47643 107541
rect 46565 107536 46612 107540
rect 46676 107538 46682 107540
rect 47526 107538 47532 107540
rect 46565 107480 46570 107536
rect 46565 107476 46612 107480
rect 46676 107478 46722 107538
rect 47486 107478 47532 107538
rect 47596 107536 47643 107540
rect 47638 107480 47643 107536
rect 46676 107476 46682 107478
rect 47526 107476 47532 107478
rect 47596 107476 47643 107480
rect 48630 107476 48636 107540
rect 48700 107538 48706 107540
rect 48773 107538 48839 107541
rect 50153 107540 50219 107541
rect 51257 107540 51323 107541
rect 52361 107540 52427 107541
rect 53465 107540 53531 107541
rect 50102 107538 50108 107540
rect 48700 107536 48839 107538
rect 48700 107480 48778 107536
rect 48834 107480 48839 107536
rect 48700 107478 48839 107480
rect 50062 107478 50108 107538
rect 50172 107536 50219 107540
rect 51206 107538 51212 107540
rect 50214 107480 50219 107536
rect 48700 107476 48706 107478
rect 46565 107475 46631 107476
rect 47577 107475 47643 107476
rect 48773 107475 48839 107478
rect 50102 107476 50108 107478
rect 50172 107476 50219 107480
rect 51166 107478 51212 107538
rect 51276 107536 51323 107540
rect 52310 107538 52316 107540
rect 51318 107480 51323 107536
rect 51206 107476 51212 107478
rect 51276 107476 51323 107480
rect 52270 107478 52316 107538
rect 52380 107536 52427 107540
rect 53414 107538 53420 107540
rect 52422 107480 52427 107536
rect 52310 107476 52316 107478
rect 52380 107476 52427 107480
rect 53374 107478 53420 107538
rect 53484 107536 53531 107540
rect 53526 107480 53531 107536
rect 53414 107476 53420 107478
rect 53484 107476 53531 107480
rect 59486 107476 59492 107540
rect 59556 107538 59562 107540
rect 59629 107538 59695 107541
rect 59556 107536 59695 107538
rect 59556 107480 59634 107536
rect 59690 107480 59695 107536
rect 59556 107478 59695 107480
rect 59556 107476 59562 107478
rect 50153 107475 50219 107476
rect 51257 107475 51323 107476
rect 52361 107475 52427 107476
rect 53465 107475 53531 107476
rect 59629 107475 59695 107478
rect 60549 107540 60615 107541
rect 61653 107540 61719 107541
rect 60549 107536 60596 107540
rect 60660 107538 60666 107540
rect 60549 107480 60554 107536
rect 60549 107476 60596 107480
rect 60660 107478 60706 107538
rect 61653 107536 61700 107540
rect 61764 107538 61770 107540
rect 62573 107538 62639 107541
rect 63585 107540 63651 107541
rect 62798 107538 62804 107540
rect 61653 107480 61658 107536
rect 60660 107476 60666 107478
rect 61653 107476 61700 107480
rect 61764 107478 61810 107538
rect 62573 107536 62804 107538
rect 62573 107480 62578 107536
rect 62634 107480 62804 107536
rect 62573 107478 62804 107480
rect 61764 107476 61770 107478
rect 60549 107475 60615 107476
rect 61653 107475 61719 107476
rect 62573 107475 62639 107478
rect 62798 107476 62804 107478
rect 62868 107476 62874 107540
rect 63534 107538 63540 107540
rect 63494 107478 63540 107538
rect 63604 107536 63651 107540
rect 63646 107480 63651 107536
rect 63534 107476 63540 107478
rect 63604 107476 63651 107480
rect 63585 107475 63651 107476
rect 63861 107540 63927 107541
rect 65149 107540 65215 107541
rect 66253 107540 66319 107541
rect 67633 107540 67699 107541
rect 63861 107536 63908 107540
rect 63972 107538 63978 107540
rect 63861 107480 63866 107536
rect 63861 107476 63908 107480
rect 63972 107478 64018 107538
rect 65149 107536 65196 107540
rect 65260 107538 65266 107540
rect 65149 107480 65154 107536
rect 63972 107476 63978 107478
rect 65149 107476 65196 107480
rect 65260 107478 65306 107538
rect 66253 107536 66300 107540
rect 66364 107538 66370 107540
rect 67582 107538 67588 107540
rect 66253 107480 66258 107536
rect 65260 107476 65266 107478
rect 66253 107476 66300 107480
rect 66364 107478 66410 107538
rect 67542 107478 67588 107538
rect 67652 107536 67699 107540
rect 67694 107480 67699 107536
rect 66364 107476 66370 107478
rect 67582 107476 67588 107478
rect 67652 107476 67699 107480
rect 63861 107475 63927 107476
rect 65149 107475 65215 107476
rect 66253 107475 66319 107476
rect 67633 107475 67699 107476
rect 68645 107540 68711 107541
rect 69749 107540 69815 107541
rect 71221 107540 71287 107541
rect 72141 107540 72207 107541
rect 73245 107540 73311 107541
rect 73705 107540 73771 107541
rect 68645 107536 68692 107540
rect 68756 107538 68762 107540
rect 68645 107480 68650 107536
rect 68645 107476 68692 107480
rect 68756 107478 68802 107538
rect 69749 107536 69796 107540
rect 69860 107538 69866 107540
rect 69749 107480 69754 107536
rect 68756 107476 68762 107478
rect 69749 107476 69796 107480
rect 69860 107478 69906 107538
rect 71221 107536 71268 107540
rect 71332 107538 71338 107540
rect 71221 107480 71226 107536
rect 69860 107476 69866 107478
rect 71221 107476 71268 107480
rect 71332 107478 71378 107538
rect 72141 107536 72188 107540
rect 72252 107538 72258 107540
rect 72141 107480 72146 107536
rect 71332 107476 71338 107478
rect 72141 107476 72188 107480
rect 72252 107478 72298 107538
rect 73245 107536 73292 107540
rect 73356 107538 73362 107540
rect 73654 107538 73660 107540
rect 73245 107480 73250 107536
rect 72252 107476 72258 107478
rect 73245 107476 73292 107480
rect 73356 107478 73402 107538
rect 73614 107478 73660 107538
rect 73724 107536 73771 107540
rect 73766 107480 73771 107536
rect 73356 107476 73362 107478
rect 73654 107476 73660 107478
rect 73724 107476 73771 107480
rect 68645 107475 68711 107476
rect 69749 107475 69815 107476
rect 71221 107475 71287 107476
rect 72141 107475 72207 107476
rect 73245 107475 73311 107476
rect 73705 107475 73771 107476
rect 74349 107540 74415 107541
rect 75637 107540 75703 107541
rect 76097 107540 76163 107541
rect 74349 107536 74396 107540
rect 74460 107538 74466 107540
rect 74349 107480 74354 107536
rect 74349 107476 74396 107480
rect 74460 107478 74506 107538
rect 75637 107536 75684 107540
rect 75748 107538 75754 107540
rect 76046 107538 76052 107540
rect 75637 107480 75642 107536
rect 74460 107476 74466 107478
rect 75637 107476 75684 107480
rect 75748 107478 75794 107538
rect 76006 107478 76052 107538
rect 76116 107536 76163 107540
rect 76158 107480 76163 107536
rect 75748 107476 75754 107478
rect 76046 107476 76052 107478
rect 76116 107476 76163 107480
rect 74349 107475 74415 107476
rect 75637 107475 75703 107476
rect 76097 107475 76163 107476
rect 77661 107538 77727 107541
rect 78489 107540 78555 107541
rect 78070 107538 78076 107540
rect 77661 107536 78076 107538
rect 77661 107480 77666 107536
rect 77722 107480 78076 107536
rect 77661 107478 78076 107480
rect 77661 107475 77727 107478
rect 78070 107476 78076 107478
rect 78140 107476 78146 107540
rect 78438 107538 78444 107540
rect 78398 107478 78444 107538
rect 78508 107536 78555 107540
rect 78550 107480 78555 107536
rect 78438 107476 78444 107478
rect 78508 107476 78555 107480
rect 78489 107475 78555 107476
rect 79133 107540 79199 107541
rect 86033 107540 86099 107541
rect 88241 107540 88307 107541
rect 93577 107540 93643 107541
rect 98545 107540 98611 107541
rect 120993 107540 121059 107541
rect 123385 107540 123451 107541
rect 79133 107536 79180 107540
rect 79244 107538 79250 107540
rect 85982 107538 85988 107540
rect 79133 107480 79138 107536
rect 79133 107476 79180 107480
rect 79244 107478 79290 107538
rect 85942 107478 85988 107538
rect 86052 107536 86099 107540
rect 88190 107538 88196 107540
rect 86094 107480 86099 107536
rect 79244 107476 79250 107478
rect 85982 107476 85988 107478
rect 86052 107476 86099 107480
rect 88150 107478 88196 107538
rect 88260 107536 88307 107540
rect 93526 107538 93532 107540
rect 88302 107480 88307 107536
rect 88190 107476 88196 107478
rect 88260 107476 88307 107480
rect 93486 107478 93532 107538
rect 93596 107536 93643 107540
rect 98494 107538 98500 107540
rect 93638 107480 93643 107536
rect 93526 107476 93532 107478
rect 93596 107476 93643 107480
rect 98454 107478 98500 107538
rect 98564 107536 98611 107540
rect 120942 107538 120948 107540
rect 98606 107480 98611 107536
rect 98494 107476 98500 107478
rect 98564 107476 98611 107480
rect 120902 107478 120948 107538
rect 121012 107536 121059 107540
rect 123334 107538 123340 107540
rect 121054 107480 121059 107536
rect 120942 107476 120948 107478
rect 121012 107476 121059 107480
rect 123294 107478 123340 107538
rect 123404 107536 123451 107540
rect 123446 107480 123451 107536
rect 123334 107476 123340 107478
rect 123404 107476 123451 107480
rect 417366 107476 417372 107540
rect 417436 107538 417442 107540
rect 418061 107538 418127 107541
rect 417436 107536 418127 107538
rect 417436 107480 418066 107536
rect 418122 107480 418127 107536
rect 417436 107478 418127 107480
rect 417436 107476 417442 107478
rect 79133 107475 79199 107476
rect 86033 107475 86099 107476
rect 88241 107475 88307 107476
rect 93577 107475 93643 107476
rect 98545 107475 98611 107476
rect 120993 107475 121059 107476
rect 123385 107475 123451 107476
rect 418061 107475 418127 107478
rect 436093 107540 436159 107541
rect 437013 107540 437079 107541
rect 438117 107540 438183 107541
rect 439589 107540 439655 107541
rect 440509 107540 440575 107541
rect 441613 107540 441679 107541
rect 443085 107540 443151 107541
rect 444189 107540 444255 107541
rect 436093 107536 436140 107540
rect 436204 107538 436210 107540
rect 436093 107480 436098 107536
rect 436093 107476 436140 107480
rect 436204 107478 436250 107538
rect 437013 107536 437060 107540
rect 437124 107538 437130 107540
rect 437013 107480 437018 107536
rect 436204 107476 436210 107478
rect 437013 107476 437060 107480
rect 437124 107478 437170 107538
rect 438117 107536 438164 107540
rect 438228 107538 438234 107540
rect 438117 107480 438122 107536
rect 437124 107476 437130 107478
rect 438117 107476 438164 107480
rect 438228 107478 438274 107538
rect 439589 107536 439636 107540
rect 439700 107538 439706 107540
rect 439589 107480 439594 107536
rect 438228 107476 438234 107478
rect 439589 107476 439636 107480
rect 439700 107478 439746 107538
rect 440509 107536 440556 107540
rect 440620 107538 440626 107540
rect 440509 107480 440514 107536
rect 439700 107476 439706 107478
rect 440509 107476 440556 107480
rect 440620 107478 440666 107538
rect 441613 107536 441660 107540
rect 441724 107538 441730 107540
rect 441613 107480 441618 107536
rect 440620 107476 440626 107478
rect 441613 107476 441660 107480
rect 441724 107478 441770 107538
rect 443085 107536 443132 107540
rect 443196 107538 443202 107540
rect 443085 107480 443090 107536
rect 441724 107476 441730 107478
rect 443085 107476 443132 107480
rect 443196 107478 443242 107538
rect 444189 107536 444236 107540
rect 444300 107538 444306 107540
rect 444189 107480 444194 107536
rect 443196 107476 443202 107478
rect 444189 107476 444236 107480
rect 444300 107478 444346 107538
rect 444300 107476 444306 107478
rect 445518 107476 445524 107540
rect 445588 107538 445594 107540
rect 445661 107538 445727 107541
rect 445588 107536 445727 107538
rect 445588 107480 445666 107536
rect 445722 107480 445727 107536
rect 445588 107478 445727 107480
rect 445588 107476 445594 107478
rect 436093 107475 436159 107476
rect 437013 107475 437079 107476
rect 438117 107475 438183 107476
rect 439589 107475 439655 107476
rect 440509 107475 440575 107476
rect 441613 107475 441679 107476
rect 443085 107475 443151 107476
rect 444189 107475 444255 107476
rect 445661 107475 445727 107478
rect 446397 107540 446463 107541
rect 446397 107536 446444 107540
rect 446508 107538 446514 107540
rect 447133 107538 447199 107541
rect 447542 107538 447548 107540
rect 446397 107480 446402 107536
rect 446397 107476 446444 107480
rect 446508 107478 446554 107538
rect 447133 107536 447548 107538
rect 447133 107480 447138 107536
rect 447194 107480 447548 107536
rect 447133 107478 447548 107480
rect 446508 107476 446514 107478
rect 446397 107475 446463 107476
rect 447133 107475 447199 107478
rect 447542 107476 447548 107478
rect 447612 107476 447618 107540
rect 448513 107538 448579 107541
rect 448646 107538 448652 107540
rect 448513 107536 448652 107538
rect 448513 107480 448518 107536
rect 448574 107480 448652 107536
rect 448513 107478 448652 107480
rect 448513 107475 448579 107478
rect 448646 107476 448652 107478
rect 448716 107476 448722 107540
rect 449893 107538 449959 107541
rect 450629 107540 450695 107541
rect 450118 107538 450124 107540
rect 449893 107536 450124 107538
rect 449893 107480 449898 107536
rect 449954 107480 450124 107536
rect 449893 107478 450124 107480
rect 449893 107475 449959 107478
rect 450118 107476 450124 107478
rect 450188 107476 450194 107540
rect 450629 107536 450676 107540
rect 450740 107538 450746 107540
rect 450629 107480 450634 107536
rect 450629 107476 450676 107480
rect 450740 107478 450786 107538
rect 450740 107476 450746 107478
rect 452326 107476 452332 107540
rect 452396 107538 452402 107540
rect 452561 107538 452627 107541
rect 452396 107536 452627 107538
rect 452396 107480 452566 107536
rect 452622 107480 452627 107536
rect 452396 107478 452627 107480
rect 452396 107476 452402 107478
rect 450629 107475 450695 107476
rect 452561 107475 452627 107478
rect 453573 107540 453639 107541
rect 454585 107540 454651 107541
rect 453573 107536 453620 107540
rect 453684 107538 453690 107540
rect 454534 107538 454540 107540
rect 453573 107480 453578 107536
rect 453573 107476 453620 107480
rect 453684 107478 453730 107538
rect 454494 107478 454540 107538
rect 454604 107536 454651 107540
rect 455781 107540 455847 107541
rect 455965 107540 456031 107541
rect 458357 107540 458423 107541
rect 459461 107540 459527 107541
rect 460657 107540 460723 107541
rect 455781 107538 455828 107540
rect 454646 107480 454651 107536
rect 453684 107476 453690 107478
rect 454534 107476 454540 107478
rect 454604 107476 454651 107480
rect 455736 107536 455828 107538
rect 455736 107480 455786 107536
rect 455736 107478 455828 107480
rect 453573 107475 453639 107476
rect 454585 107475 454651 107476
rect 455781 107476 455828 107478
rect 455892 107476 455898 107540
rect 455965 107536 456012 107540
rect 456076 107538 456082 107540
rect 455965 107480 455970 107536
rect 455965 107476 456012 107480
rect 456076 107478 456122 107538
rect 458357 107536 458404 107540
rect 458468 107538 458474 107540
rect 458357 107480 458362 107536
rect 456076 107476 456082 107478
rect 458357 107476 458404 107480
rect 458468 107478 458514 107538
rect 459461 107536 459508 107540
rect 459572 107538 459578 107540
rect 460606 107538 460612 107540
rect 459461 107480 459466 107536
rect 458468 107476 458474 107478
rect 459461 107476 459508 107480
rect 459572 107478 459618 107538
rect 460566 107478 460612 107538
rect 460676 107536 460723 107540
rect 460718 107480 460723 107536
rect 459572 107476 459578 107478
rect 460606 107476 460612 107478
rect 460676 107476 460723 107480
rect 455781 107475 455847 107476
rect 455965 107475 456031 107476
rect 458357 107475 458423 107476
rect 459461 107475 459527 107476
rect 460657 107475 460723 107476
rect 461669 107540 461735 107541
rect 462773 107540 462839 107541
rect 463877 107540 463943 107541
rect 465165 107540 465231 107541
rect 461669 107536 461716 107540
rect 461780 107538 461786 107540
rect 461669 107480 461674 107536
rect 461669 107476 461716 107480
rect 461780 107478 461826 107538
rect 462773 107536 462820 107540
rect 462884 107538 462890 107540
rect 462773 107480 462778 107536
rect 461780 107476 461786 107478
rect 462773 107476 462820 107480
rect 462884 107478 462930 107538
rect 463877 107536 463924 107540
rect 463988 107538 463994 107540
rect 463877 107480 463882 107536
rect 462884 107476 462890 107478
rect 463877 107476 463924 107480
rect 463988 107478 464034 107538
rect 465165 107536 465212 107540
rect 465276 107538 465282 107540
rect 465717 107538 465783 107541
rect 466310 107538 466316 107540
rect 465165 107480 465170 107536
rect 463988 107476 463994 107478
rect 465165 107476 465212 107480
rect 465276 107478 465322 107538
rect 465717 107536 466316 107538
rect 465717 107480 465722 107536
rect 465778 107480 466316 107536
rect 465717 107478 466316 107480
rect 465276 107476 465282 107478
rect 461669 107475 461735 107476
rect 462773 107475 462839 107476
rect 463877 107475 463943 107476
rect 465165 107475 465231 107476
rect 465717 107475 465783 107478
rect 466310 107476 466316 107478
rect 466380 107476 466386 107540
rect 467005 107538 467071 107541
rect 468661 107540 468727 107541
rect 469765 107540 469831 107541
rect 467598 107538 467604 107540
rect 467005 107536 467604 107538
rect 467005 107480 467010 107536
rect 467066 107480 467604 107536
rect 467005 107478 467604 107480
rect 467005 107475 467071 107478
rect 467598 107476 467604 107478
rect 467668 107476 467674 107540
rect 468661 107536 468708 107540
rect 468772 107538 468778 107540
rect 468661 107480 468666 107536
rect 468661 107476 468708 107480
rect 468772 107478 468818 107538
rect 469765 107536 469812 107540
rect 469876 107538 469882 107540
rect 471145 107538 471211 107541
rect 471278 107538 471284 107540
rect 469765 107480 469770 107536
rect 468772 107476 468778 107478
rect 469765 107476 469812 107480
rect 469876 107478 469922 107538
rect 471145 107536 471284 107538
rect 471145 107480 471150 107536
rect 471206 107480 471284 107536
rect 471145 107478 471284 107480
rect 469876 107476 469882 107478
rect 468661 107475 468727 107476
rect 469765 107475 469831 107476
rect 471145 107475 471211 107478
rect 471278 107476 471284 107478
rect 471348 107476 471354 107540
rect 472065 107538 472131 107541
rect 473353 107540 473419 107541
rect 472198 107538 472204 107540
rect 472065 107536 472204 107538
rect 472065 107480 472070 107536
rect 472126 107480 472204 107536
rect 472065 107478 472204 107480
rect 472065 107475 472131 107478
rect 472198 107476 472204 107478
rect 472268 107476 472274 107540
rect 473302 107538 473308 107540
rect 473262 107478 473308 107538
rect 473372 107536 473419 107540
rect 473414 107480 473419 107536
rect 473302 107476 473308 107478
rect 473372 107476 473419 107480
rect 473353 107475 473419 107476
rect 474365 107540 474431 107541
rect 475653 107540 475719 107541
rect 478045 107540 478111 107541
rect 479149 107540 479215 107541
rect 474365 107536 474412 107540
rect 474476 107538 474482 107540
rect 474365 107480 474370 107536
rect 474365 107476 474412 107480
rect 474476 107478 474522 107538
rect 475653 107536 475700 107540
rect 475764 107538 475770 107540
rect 475653 107480 475658 107536
rect 474476 107476 474482 107478
rect 475653 107476 475700 107480
rect 475764 107478 475810 107538
rect 478045 107536 478092 107540
rect 478156 107538 478162 107540
rect 478045 107480 478050 107536
rect 475764 107476 475770 107478
rect 478045 107476 478092 107480
rect 478156 107478 478202 107538
rect 479149 107536 479196 107540
rect 479260 107538 479266 107540
rect 479149 107480 479154 107536
rect 478156 107476 478162 107478
rect 479149 107476 479196 107480
rect 479260 107478 479306 107538
rect 479260 107476 479266 107478
rect 474365 107475 474431 107476
rect 475653 107475 475719 107476
rect 478045 107475 478111 107476
rect 479149 107475 479215 107476
rect 19006 107340 19012 107404
rect 19076 107402 19082 107404
rect 41822 107402 41828 107404
rect 19076 107342 41828 107402
rect 19076 107340 19082 107342
rect 41822 107340 41828 107342
rect 41892 107340 41898 107404
rect 57094 107340 57100 107404
rect 57164 107402 57170 107404
rect 61745 107402 61811 107405
rect 57164 107400 61811 107402
rect 57164 107344 61750 107400
rect 61806 107344 61811 107400
rect 57164 107342 61811 107344
rect 57164 107340 57170 107342
rect 61745 107339 61811 107342
rect 70894 107340 70900 107404
rect 70964 107402 70970 107404
rect 191230 107402 191236 107404
rect 70964 107342 191236 107402
rect 70964 107340 70970 107342
rect 191230 107340 191236 107342
rect 191300 107340 191306 107404
rect 388713 107402 388779 107405
rect 463550 107402 463556 107404
rect 388713 107400 463556 107402
rect 388713 107344 388718 107400
rect 388774 107344 463556 107400
rect 388713 107342 463556 107344
rect 388713 107339 388779 107342
rect 463550 107340 463556 107342
rect 463620 107340 463626 107404
rect 18413 107266 18479 107269
rect 58014 107266 58020 107268
rect 18413 107264 58020 107266
rect 18413 107208 18418 107264
rect 18474 107208 58020 107264
rect 18413 107206 58020 107208
rect 18413 107203 18479 107206
rect 58014 107204 58020 107206
rect 58084 107266 58090 107268
rect 76966 107266 76972 107268
rect 58084 107206 76972 107266
rect 58084 107204 58090 107206
rect 76966 107204 76972 107206
rect 77036 107204 77042 107268
rect 81014 107204 81020 107268
rect 81084 107266 81090 107268
rect 187366 107266 187372 107268
rect 81084 107206 187372 107266
rect 81084 107204 81090 107206
rect 187366 107204 187372 107206
rect 187436 107204 187442 107268
rect 418797 107266 418863 107269
rect 478454 107266 478460 107268
rect 418797 107264 478460 107266
rect 418797 107208 418802 107264
rect 418858 107208 478460 107264
rect 418797 107206 478460 107208
rect 418797 107203 418863 107206
rect 478454 107204 478460 107206
rect 478524 107204 478530 107268
rect 54518 107068 54524 107132
rect 54588 107130 54594 107132
rect 55121 107130 55187 107133
rect 54588 107128 55187 107130
rect 54588 107072 55126 107128
rect 55182 107072 55187 107128
rect 54588 107070 55187 107072
rect 54588 107068 54594 107070
rect 55121 107067 55187 107070
rect 55765 107132 55831 107133
rect 55765 107128 55812 107132
rect 55876 107130 55882 107132
rect 55765 107072 55770 107128
rect 55765 107068 55812 107072
rect 55876 107070 55922 107130
rect 55876 107068 55882 107070
rect 83590 107068 83596 107132
rect 83660 107130 83666 107132
rect 186998 107130 187004 107132
rect 83660 107070 187004 107130
rect 83660 107068 83666 107070
rect 186998 107068 187004 107070
rect 187068 107068 187074 107132
rect 390093 107130 390159 107133
rect 448278 107130 448284 107132
rect 390093 107128 448284 107130
rect 390093 107072 390098 107128
rect 390154 107072 448284 107128
rect 390093 107070 448284 107072
rect 55765 107067 55831 107068
rect 390093 107067 390159 107070
rect 448278 107068 448284 107070
rect 448348 107068 448354 107132
rect 453430 107068 453436 107132
rect 453500 107130 453506 107132
rect 453941 107130 454007 107133
rect 453500 107128 454007 107130
rect 453500 107072 453946 107128
rect 454002 107072 454007 107128
rect 453500 107070 454007 107072
rect 453500 107068 453506 107070
rect 453941 107067 454007 107070
rect 457989 107130 458055 107133
rect 476982 107130 476988 107132
rect 457989 107128 476988 107130
rect 457989 107072 457994 107128
rect 458050 107072 476988 107128
rect 457989 107070 476988 107072
rect 457989 107067 458055 107070
rect 476982 107068 476988 107070
rect 477052 107068 477058 107132
rect 103462 106932 103468 106996
rect 103532 106994 103538 106996
rect 191414 106994 191420 106996
rect 103532 106934 191420 106994
rect 103532 106932 103538 106934
rect 191414 106932 191420 106934
rect 191484 106932 191490 106996
rect 419022 106932 419028 106996
rect 419092 106994 419098 106996
rect 473486 106994 473492 106996
rect 419092 106934 473492 106994
rect 419092 106932 419098 106934
rect 473486 106932 473492 106934
rect 473556 106932 473562 106996
rect 115790 106796 115796 106860
rect 115860 106858 115866 106860
rect 184054 106858 184060 106860
rect 115860 106798 184060 106858
rect 115860 106796 115866 106798
rect 184054 106796 184060 106798
rect 184124 106796 184130 106860
rect 58566 106660 58572 106724
rect 58636 106722 58642 106724
rect 182081 106722 182147 106725
rect 58636 106720 182147 106722
rect 58636 106664 182086 106720
rect 182142 106664 182147 106720
rect 58636 106662 182147 106664
rect 58636 106660 58642 106662
rect 182081 106659 182147 106662
rect 388529 106722 388595 106725
rect 511022 106722 511028 106724
rect 388529 106720 511028 106722
rect 388529 106664 388534 106720
rect 388590 106664 511028 106720
rect 388529 106662 511028 106664
rect 388529 106659 388595 106662
rect 511022 106660 511028 106662
rect 511092 106660 511098 106724
rect 57053 106316 57119 106317
rect 57053 106312 57100 106316
rect 57164 106314 57170 106316
rect 57053 106256 57058 106312
rect 57053 106252 57100 106256
rect 57164 106254 57210 106314
rect 57164 106252 57170 106254
rect 57053 106251 57119 106252
rect 350942 106116 350948 106180
rect 351012 106178 351018 106180
rect 351177 106178 351243 106181
rect 351012 106176 351243 106178
rect 351012 106120 351182 106176
rect 351238 106120 351243 106176
rect 351012 106118 351243 106120
rect 351012 106116 351018 106118
rect 351177 106115 351243 106118
rect 191598 105708 191604 105772
rect 191668 105770 191674 105772
rect 580901 105770 580967 105773
rect 191668 105768 580967 105770
rect 191668 105712 580906 105768
rect 580962 105712 580967 105768
rect 191668 105710 580967 105712
rect 191668 105708 191674 105710
rect 580901 105707 580967 105710
rect 188838 105572 188844 105636
rect 188908 105634 188914 105636
rect 580441 105634 580507 105637
rect 188908 105632 580507 105634
rect 188908 105576 580446 105632
rect 580502 105576 580507 105632
rect 188908 105574 580507 105576
rect 188908 105572 188914 105574
rect 580441 105571 580507 105574
rect 188654 105436 188660 105500
rect 188724 105498 188730 105500
rect 580717 105498 580783 105501
rect 188724 105496 580783 105498
rect 188724 105440 580722 105496
rect 580778 105440 580783 105496
rect 188724 105438 580783 105440
rect 188724 105436 188730 105438
rect 580717 105435 580783 105438
rect 150801 105364 150867 105365
rect 150750 105362 150756 105364
rect 150710 105302 150756 105362
rect 150820 105360 150867 105364
rect 150862 105304 150867 105360
rect 150750 105300 150756 105302
rect 150820 105300 150867 105304
rect 150801 105299 150867 105300
rect 550725 105364 550791 105365
rect 550725 105360 550772 105364
rect 550836 105362 550842 105364
rect 550725 105304 550730 105360
rect 550725 105300 550772 105304
rect 550836 105302 550882 105362
rect 550836 105300 550842 105302
rect 550725 105299 550791 105300
rect 580349 99514 580415 99517
rect 583520 99514 584960 99604
rect 580349 99512 584960 99514
rect 580349 99456 580354 99512
rect 580410 99456 584960 99512
rect 580349 99454 584960 99456
rect 580349 99451 580415 99454
rect 558913 99378 558979 99381
rect 556570 99376 558979 99378
rect 556570 99320 558918 99376
rect 558974 99320 558979 99376
rect 583520 99364 584960 99454
rect 556570 99318 558979 99320
rect 158713 99242 158779 99245
rect 158897 99242 158963 99245
rect 359733 99242 359799 99245
rect 360101 99242 360167 99245
rect 156558 99240 158963 99242
rect 156558 99184 158718 99240
rect 158774 99184 158902 99240
rect 158958 99184 158963 99240
rect 156558 99182 158963 99184
rect 356562 99240 360167 99242
rect 356562 99184 359738 99240
rect 359794 99184 360106 99240
rect 360162 99184 360167 99240
rect 556570 99190 556630 99318
rect 558913 99315 558979 99318
rect 356562 99182 360167 99184
rect 158713 99179 158779 99182
rect 158897 99179 158963 99182
rect 359733 99179 359799 99182
rect 360101 99179 360167 99182
rect -960 97610 480 97700
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 18454 96658 18460 96660
rect 6870 96598 18460 96658
rect 18454 96596 18460 96598
rect 18524 96596 18530 96660
rect 580901 86186 580967 86189
rect 583520 86186 584960 86276
rect 580901 86184 584960 86186
rect 580901 86128 580906 86184
rect 580962 86128 584960 86184
rect 580901 86126 584960 86128
rect 580901 86123 580967 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3693 84690 3759 84693
rect -960 84688 3759 84690
rect -960 84632 3698 84688
rect 3754 84632 3759 84688
rect -960 84630 3759 84632
rect -960 84540 480 84630
rect 3693 84627 3759 84630
rect 580717 72994 580783 72997
rect 583520 72994 584960 73084
rect 580717 72992 584960 72994
rect 580717 72936 580722 72992
rect 580778 72936 584960 72992
rect 580717 72934 584960 72936
rect 580717 72931 580783 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 580441 59666 580507 59669
rect 583520 59666 584960 59756
rect 580441 59664 584960 59666
rect 580441 59608 580446 59664
rect 580502 59608 584960 59664
rect 580441 59606 584960 59608
rect 580441 59603 580507 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 17309 56946 17375 56949
rect 216673 56946 216739 56949
rect 417325 56946 417391 56949
rect 17309 56944 19442 56946
rect 17309 56888 17314 56944
rect 17370 56924 19442 56944
rect 216673 56944 219450 56946
rect 17370 56888 20056 56924
rect 17309 56886 20056 56888
rect 17309 56883 17375 56886
rect 19382 56864 20056 56886
rect 216673 56888 216678 56944
rect 216734 56924 219450 56944
rect 417325 56944 419458 56946
rect 216734 56888 220064 56924
rect 216673 56886 220064 56888
rect 216673 56883 216739 56886
rect 219390 56864 220064 56886
rect 417325 56888 417330 56944
rect 417386 56924 419458 56944
rect 417386 56888 420072 56924
rect 417325 56886 420072 56888
rect 417325 56883 417391 56886
rect 419398 56864 420072 56886
rect 17401 55994 17467 55997
rect 216673 55994 216739 55997
rect 17401 55992 19442 55994
rect 17401 55936 17406 55992
rect 17462 55972 19442 55992
rect 216673 55992 219450 55994
rect 17462 55936 20056 55972
rect 17401 55934 20056 55936
rect 17401 55931 17467 55934
rect 19382 55912 20056 55934
rect 216673 55936 216678 55992
rect 216734 55972 219450 55992
rect 216734 55936 220064 55972
rect 216673 55934 220064 55936
rect 216673 55931 216739 55934
rect 219390 55912 220064 55934
rect 417182 55932 417188 55996
rect 417252 55994 417258 55996
rect 417252 55972 419458 55994
rect 417252 55934 420072 55972
rect 417252 55932 417258 55934
rect 419398 55912 420072 55934
rect 17677 53818 17743 53821
rect 216673 53818 216739 53821
rect 417601 53818 417667 53821
rect 17677 53816 19442 53818
rect 17677 53760 17682 53816
rect 17738 53796 19442 53816
rect 216673 53816 219450 53818
rect 17738 53760 20056 53796
rect 17677 53758 20056 53760
rect 17677 53755 17743 53758
rect 19382 53736 20056 53758
rect 216673 53760 216678 53816
rect 216734 53796 219450 53816
rect 417601 53816 419458 53818
rect 216734 53760 220064 53796
rect 216673 53758 220064 53760
rect 216673 53755 216739 53758
rect 219390 53736 220064 53758
rect 417601 53760 417606 53816
rect 417662 53796 419458 53816
rect 417662 53760 420072 53796
rect 417601 53758 420072 53760
rect 417601 53755 417667 53758
rect 419398 53736 420072 53758
rect 17493 52866 17559 52869
rect 216765 52866 216831 52869
rect 17493 52864 19442 52866
rect 17493 52808 17498 52864
rect 17554 52844 19442 52864
rect 216765 52864 219450 52866
rect 17554 52808 20056 52844
rect 17493 52806 20056 52808
rect 17493 52803 17559 52806
rect 19382 52784 20056 52806
rect 216765 52808 216770 52864
rect 216826 52844 219450 52864
rect 216826 52808 220064 52844
rect 216765 52806 220064 52808
rect 216765 52803 216831 52806
rect 219390 52784 220064 52806
rect 417734 52804 417740 52868
rect 417804 52866 417810 52868
rect 417804 52844 419458 52866
rect 417804 52806 420072 52844
rect 417804 52804 417810 52806
rect 419398 52784 420072 52806
rect 17769 51098 17835 51101
rect 216765 51098 216831 51101
rect 417509 51098 417575 51101
rect 17769 51096 19810 51098
rect 17769 51040 17774 51096
rect 17830 51076 19810 51096
rect 216765 51096 220002 51098
rect 17830 51040 20056 51076
rect 17769 51038 20056 51040
rect 17769 51035 17835 51038
rect 19750 51016 20056 51038
rect 216765 51040 216770 51096
rect 216826 51076 220002 51096
rect 417509 51096 420010 51098
rect 216826 51040 220064 51076
rect 216765 51038 220064 51040
rect 216765 51035 216831 51038
rect 219942 51016 220064 51038
rect 417509 51040 417514 51096
rect 417570 51076 420010 51096
rect 417570 51040 420072 51076
rect 417509 51038 420072 51040
rect 417509 51035 417575 51038
rect 419950 51016 420072 51038
rect 17585 50010 17651 50013
rect 216673 50010 216739 50013
rect 417233 50010 417299 50013
rect 17585 50008 19442 50010
rect 17585 49952 17590 50008
rect 17646 49988 19442 50008
rect 216673 50008 219450 50010
rect 17646 49952 20056 49988
rect 17585 49950 20056 49952
rect 17585 49947 17651 49950
rect 19382 49928 20056 49950
rect 216673 49952 216678 50008
rect 216734 49988 219450 50008
rect 417233 50008 419458 50010
rect 216734 49952 220064 49988
rect 216673 49950 220064 49952
rect 216673 49947 216739 49950
rect 219390 49928 220064 49950
rect 417233 49952 417238 50008
rect 417294 49988 419458 50008
rect 417294 49952 420072 49988
rect 417233 49950 420072 49952
rect 417233 49947 417299 49950
rect 419398 49928 420072 49950
rect 17861 48242 17927 48245
rect 216673 48242 216739 48245
rect 17861 48240 19442 48242
rect 17861 48184 17866 48240
rect 17922 48220 19442 48240
rect 216673 48240 219450 48242
rect 17922 48184 20056 48220
rect 17861 48182 20056 48184
rect 17861 48179 17927 48182
rect 19382 48160 20056 48182
rect 216673 48184 216678 48240
rect 216734 48220 219450 48240
rect 216734 48184 220064 48220
rect 216673 48182 220064 48184
rect 216673 48179 216739 48182
rect 219390 48160 220064 48182
rect 417918 48180 417924 48244
rect 417988 48242 417994 48244
rect 417988 48220 419458 48242
rect 417988 48182 420072 48220
rect 417988 48180 417994 48182
rect 419398 48160 420072 48182
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3325 45522 3391 45525
rect -960 45520 3391 45522
rect -960 45464 3330 45520
rect 3386 45464 3391 45520
rect -960 45462 3391 45464
rect -960 45372 480 45462
rect 3325 45459 3391 45462
rect 580809 33146 580875 33149
rect 583520 33146 584960 33236
rect 580809 33144 584960 33146
rect 580809 33088 580814 33144
rect 580870 33088 584960 33144
rect 580809 33086 584960 33088
rect 580809 33083 580875 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3325 32466 3391 32469
rect -960 32464 3391 32466
rect -960 32408 3330 32464
rect 3386 32408 3391 32464
rect -960 32406 3391 32408
rect -960 32316 480 32406
rect 3325 32403 3391 32406
rect 17033 30018 17099 30021
rect 17033 30016 19442 30018
rect 17033 29960 17038 30016
rect 17094 29996 19442 30016
rect 17094 29960 20056 29996
rect 17033 29958 20056 29960
rect 17033 29955 17099 29958
rect 19382 29936 20056 29958
rect 190310 29956 190316 30020
rect 190380 30018 190386 30020
rect 417417 30018 417483 30021
rect 190380 29996 219450 30018
rect 417417 30016 419458 30018
rect 190380 29958 220064 29996
rect 190380 29956 190386 29958
rect 219390 29936 220064 29958
rect 417417 29960 417422 30016
rect 417478 29996 419458 30016
rect 417478 29960 420072 29996
rect 417417 29958 420072 29960
rect 417417 29955 417483 29958
rect 419398 29936 420072 29958
rect 217317 28522 217383 28525
rect 217182 28520 217383 28522
rect 217182 28464 217322 28520
rect 217378 28464 217383 28520
rect 217182 28462 217383 28464
rect 17217 28386 17283 28389
rect 17217 28384 19442 28386
rect 17217 28328 17222 28384
rect 17278 28364 19442 28384
rect 17278 28328 20056 28364
rect 17217 28326 20056 28328
rect 17217 28323 17283 28326
rect 19382 28304 20056 28326
rect 19190 28052 19196 28116
rect 19260 28114 19266 28116
rect 217182 28114 217242 28462
rect 217317 28459 217383 28462
rect 217317 28386 217383 28389
rect 416865 28386 416931 28389
rect 417785 28386 417851 28389
rect 217317 28384 219450 28386
rect 217317 28328 217322 28384
rect 217378 28364 219450 28384
rect 416865 28384 419458 28386
rect 217378 28328 220064 28364
rect 217317 28326 220064 28328
rect 217317 28323 217383 28326
rect 219390 28304 220064 28326
rect 416865 28328 416870 28384
rect 416926 28328 417790 28384
rect 417846 28364 419458 28384
rect 417846 28328 420072 28364
rect 416865 28326 420072 28328
rect 416865 28323 416931 28326
rect 417785 28323 417851 28326
rect 419398 28304 420072 28326
rect 416773 28114 416839 28117
rect 19260 28092 19810 28114
rect 217182 28092 219450 28114
rect 416773 28112 419458 28114
rect 19260 28054 20056 28092
rect 217182 28054 220064 28092
rect 19260 28052 19266 28054
rect 19750 28032 20056 28054
rect 219390 28032 220064 28054
rect 416773 28056 416778 28112
rect 416834 28092 419458 28112
rect 416834 28056 420072 28092
rect 416773 28054 420072 28056
rect 416773 28051 416839 28054
rect 419398 28032 420072 28054
rect 460657 19820 460723 19821
rect 488257 19820 488323 19821
rect 460657 19816 460670 19820
rect 460734 19818 460740 19820
rect 488257 19818 488278 19820
rect 460657 19760 460662 19816
rect 460657 19756 460670 19760
rect 460734 19758 460814 19818
rect 488186 19816 488278 19818
rect 488186 19760 488262 19816
rect 488186 19758 488278 19760
rect 460734 19756 460740 19758
rect 488257 19756 488278 19758
rect 488342 19756 488348 19820
rect 580625 19818 580691 19821
rect 583520 19818 584960 19908
rect 580625 19816 584960 19818
rect 580625 19760 580630 19816
rect 580686 19760 584960 19816
rect 580625 19758 584960 19760
rect 460657 19755 460723 19756
rect 488257 19755 488323 19756
rect 580625 19755 580691 19758
rect 447593 19684 447659 19685
rect 448697 19684 448763 19685
rect 450077 19684 450143 19685
rect 455965 19684 456031 19685
rect 473353 19684 473419 19685
rect 491017 19684 491083 19685
rect 447593 19680 447614 19684
rect 447678 19682 447684 19684
rect 447593 19624 447598 19680
rect 447593 19620 447614 19624
rect 447678 19622 447750 19682
rect 447678 19620 447684 19622
rect 448696 19620 448702 19684
rect 448766 19682 448772 19684
rect 450056 19682 450062 19684
rect 448766 19622 448854 19682
rect 449986 19622 450062 19682
rect 450126 19680 450143 19684
rect 455904 19682 455910 19684
rect 450138 19624 450143 19680
rect 448766 19620 448772 19622
rect 450056 19620 450062 19622
rect 450126 19620 450143 19624
rect 455874 19622 455910 19682
rect 455974 19680 456031 19684
rect 456026 19624 456031 19680
rect 455904 19620 455910 19622
rect 455974 19620 456031 19624
rect 473312 19620 473318 19684
rect 473382 19682 473419 19684
rect 473382 19680 473474 19682
rect 473414 19624 473474 19680
rect 473382 19622 473474 19624
rect 473382 19620 473419 19622
rect 490992 19620 490998 19684
rect 491062 19682 491083 19684
rect 493409 19684 493475 19685
rect 493409 19682 493446 19684
rect 491062 19680 491154 19682
rect 491078 19624 491154 19680
rect 491062 19622 491154 19624
rect 493354 19680 493446 19682
rect 493354 19624 493414 19680
rect 493354 19622 493446 19624
rect 491062 19620 491083 19622
rect 447593 19619 447659 19620
rect 448697 19619 448763 19620
rect 450077 19619 450143 19620
rect 455965 19619 456031 19620
rect 473353 19619 473419 19620
rect 491017 19619 491083 19620
rect 493409 19620 493446 19622
rect 493510 19620 493516 19684
rect 583520 19668 584960 19758
rect 493409 19619 493475 19620
rect 52361 19548 52427 19549
rect 53465 19548 53531 19549
rect 55949 19548 56015 19549
rect 52361 19544 52374 19548
rect 52438 19546 52444 19548
rect 53456 19546 53462 19548
rect -960 19410 480 19500
rect 52361 19488 52366 19544
rect 52361 19484 52374 19488
rect 52438 19486 52518 19546
rect 53374 19486 53462 19546
rect 52438 19484 52444 19486
rect 53456 19484 53462 19486
rect 53526 19484 53532 19548
rect 55904 19546 55910 19548
rect 55858 19486 55910 19546
rect 55974 19544 56015 19548
rect 285949 19548 286015 19549
rect 285949 19546 285966 19548
rect 56010 19488 56015 19544
rect 55904 19484 55910 19486
rect 55974 19484 56015 19488
rect 285874 19544 285966 19546
rect 285874 19488 285954 19544
rect 285874 19486 285966 19488
rect 52361 19483 52427 19484
rect 53465 19483 53531 19484
rect 55949 19483 56015 19484
rect 285949 19484 285966 19486
rect 286030 19484 286036 19548
rect 402329 19546 402395 19549
rect 468293 19548 468359 19549
rect 495893 19548 495959 19549
rect 500953 19548 501019 19549
rect 503529 19548 503595 19549
rect 461072 19546 461078 19548
rect 402329 19544 461078 19546
rect 402329 19488 402334 19544
rect 402390 19488 461078 19544
rect 402329 19486 461078 19488
rect 285949 19483 286015 19484
rect 402329 19483 402395 19486
rect 461072 19484 461078 19486
rect 461142 19484 461148 19548
rect 468280 19484 468286 19548
rect 468350 19546 468359 19548
rect 485960 19546 485966 19548
rect 468350 19544 468442 19546
rect 468354 19488 468442 19544
rect 468350 19486 468442 19488
rect 470550 19486 485966 19546
rect 468350 19484 468359 19486
rect 468293 19483 468359 19484
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 405365 19410 405431 19413
rect 470550 19410 470610 19486
rect 485960 19484 485966 19486
rect 486030 19484 486036 19548
rect 495888 19546 495894 19548
rect 495802 19486 495894 19546
rect 495888 19484 495894 19486
rect 495958 19484 495964 19548
rect 500920 19484 500926 19548
rect 500990 19546 501019 19548
rect 500990 19544 501082 19546
rect 501014 19488 501082 19544
rect 500990 19486 501082 19488
rect 500990 19484 501019 19486
rect 503504 19484 503510 19548
rect 503574 19546 503595 19548
rect 503574 19544 503666 19546
rect 503590 19488 503666 19544
rect 503574 19486 503666 19488
rect 503574 19484 503595 19486
rect 495893 19483 495959 19484
rect 500953 19483 501019 19484
rect 503529 19483 503595 19484
rect 405365 19408 470610 19410
rect 405365 19352 405370 19408
rect 405426 19352 470610 19408
rect 405365 19350 470610 19352
rect 405365 19347 405431 19350
rect 95969 19276 96035 19277
rect 100937 19276 101003 19277
rect 103697 19276 103763 19277
rect 95918 19212 95924 19276
rect 95988 19274 96035 19276
rect 95988 19272 96080 19274
rect 96030 19216 96080 19272
rect 95988 19214 96080 19216
rect 95988 19212 96035 19214
rect 100886 19212 100892 19276
rect 100956 19274 101003 19276
rect 100956 19272 101048 19274
rect 100998 19216 101048 19272
rect 100956 19214 101048 19216
rect 100956 19212 101003 19214
rect 103646 19212 103652 19276
rect 103716 19274 103763 19276
rect 103716 19272 103808 19274
rect 103758 19216 103808 19272
rect 103716 19214 103808 19216
rect 103716 19212 103763 19214
rect 118550 19212 118556 19276
rect 118620 19274 118626 19276
rect 173709 19274 173775 19277
rect 244273 19276 244339 19277
rect 118620 19272 173775 19274
rect 118620 19216 173714 19272
rect 173770 19216 173775 19272
rect 118620 19214 173775 19216
rect 118620 19212 118626 19214
rect 95969 19211 96035 19212
rect 100937 19211 101003 19212
rect 103697 19211 103763 19212
rect 173709 19211 173775 19214
rect 185158 19212 185164 19276
rect 185228 19274 185234 19276
rect 240542 19274 240548 19276
rect 185228 19214 240548 19274
rect 185228 19212 185234 19214
rect 240542 19212 240548 19214
rect 240612 19212 240618 19276
rect 244222 19212 244228 19276
rect 244292 19274 244339 19276
rect 245285 19276 245351 19277
rect 246389 19276 246455 19277
rect 245285 19274 245332 19276
rect 244292 19272 244384 19274
rect 244334 19216 244384 19272
rect 244292 19214 244384 19216
rect 245240 19272 245332 19274
rect 245240 19216 245290 19272
rect 245240 19214 245332 19216
rect 244292 19212 244339 19214
rect 244273 19211 244339 19212
rect 245285 19212 245332 19214
rect 245396 19212 245402 19276
rect 246389 19274 246436 19276
rect 246344 19272 246436 19274
rect 246344 19216 246394 19272
rect 246344 19214 246436 19216
rect 246389 19212 246436 19214
rect 246500 19212 246506 19276
rect 415894 19212 415900 19276
rect 415964 19274 415970 19276
rect 485037 19274 485103 19277
rect 498469 19276 498535 19277
rect 498469 19274 498516 19276
rect 415964 19272 485103 19274
rect 415964 19216 485042 19272
rect 485098 19216 485103 19272
rect 415964 19214 485103 19216
rect 498424 19272 498516 19274
rect 498424 19216 498474 19272
rect 498424 19214 498516 19216
rect 415964 19212 415970 19214
rect 245285 19211 245351 19212
rect 246389 19211 246455 19212
rect 485037 19211 485103 19214
rect 498469 19212 498516 19214
rect 498580 19212 498586 19276
rect 501045 19274 501111 19277
rect 520958 19274 520964 19276
rect 501045 19272 520964 19274
rect 501045 19216 501050 19272
rect 501106 19216 520964 19272
rect 501045 19214 520964 19216
rect 498469 19211 498535 19212
rect 501045 19211 501111 19214
rect 520958 19212 520964 19214
rect 521028 19212 521034 19276
rect 86033 19140 86099 19141
rect 91001 19140 91067 19141
rect 85982 19076 85988 19140
rect 86052 19138 86099 19140
rect 86052 19136 86144 19138
rect 86094 19080 86144 19136
rect 86052 19078 86144 19080
rect 86052 19076 86099 19078
rect 90950 19076 90956 19140
rect 91020 19138 91067 19140
rect 91020 19136 91112 19138
rect 91062 19080 91112 19136
rect 91020 19078 91112 19080
rect 91020 19076 91067 19078
rect 120942 19076 120948 19140
rect 121012 19138 121018 19140
rect 173525 19138 173591 19141
rect 121012 19136 173591 19138
rect 121012 19080 173530 19136
rect 173586 19080 173591 19136
rect 121012 19078 173591 19080
rect 121012 19076 121018 19078
rect 86033 19075 86099 19076
rect 91001 19075 91067 19076
rect 173525 19075 173591 19078
rect 185577 19138 185643 19141
rect 248229 19140 248295 19141
rect 250069 19140 250135 19141
rect 239622 19138 239628 19140
rect 185577 19136 239628 19138
rect 185577 19080 185582 19136
rect 185638 19080 239628 19136
rect 185577 19078 239628 19080
rect 185577 19075 185643 19078
rect 239622 19076 239628 19078
rect 239692 19076 239698 19140
rect 248229 19138 248276 19140
rect 248184 19136 248276 19138
rect 248184 19080 248234 19136
rect 248184 19078 248276 19080
rect 248229 19076 248276 19078
rect 248340 19076 248346 19140
rect 250069 19138 250116 19140
rect 250024 19136 250116 19138
rect 250024 19080 250074 19136
rect 250024 19078 250116 19080
rect 250069 19076 250116 19078
rect 250180 19076 250186 19140
rect 418102 19076 418108 19140
rect 418172 19138 418178 19140
rect 418429 19138 418495 19141
rect 418172 19136 418495 19138
rect 418172 19080 418434 19136
rect 418490 19080 418495 19136
rect 418172 19078 418495 19080
rect 418172 19076 418178 19078
rect 248229 19075 248295 19076
rect 250069 19075 250135 19076
rect 418429 19075 418495 19078
rect 418838 19076 418844 19140
rect 418908 19138 418914 19140
rect 518382 19138 518388 19140
rect 418908 19078 518388 19138
rect 418908 19076 418914 19078
rect 518382 19076 518388 19078
rect 518452 19076 518458 19140
rect 76097 19004 76163 19005
rect 81065 19004 81131 19005
rect 76046 18940 76052 19004
rect 76116 19002 76163 19004
rect 76116 19000 76208 19002
rect 76158 18944 76208 19000
rect 76116 18942 76208 18944
rect 76116 18940 76163 18942
rect 81014 18940 81020 19004
rect 81084 19002 81131 19004
rect 188337 19002 188403 19005
rect 247493 19004 247559 19005
rect 250621 19004 250687 19005
rect 515765 19004 515831 19005
rect 241646 19002 241652 19004
rect 81084 19000 81176 19002
rect 81126 18944 81176 19000
rect 81084 18942 81176 18944
rect 188337 19000 241652 19002
rect 188337 18944 188342 19000
rect 188398 18944 241652 19000
rect 188337 18942 241652 18944
rect 81084 18940 81131 18942
rect 76097 18939 76163 18940
rect 81065 18939 81131 18940
rect 188337 18939 188403 18942
rect 241646 18940 241652 18942
rect 241716 18940 241722 19004
rect 247493 19002 247540 19004
rect 247448 19000 247540 19002
rect 247448 18944 247498 19000
rect 247448 18942 247540 18944
rect 247493 18940 247540 18942
rect 247604 18940 247610 19004
rect 250621 19002 250668 19004
rect 250576 19000 250668 19002
rect 250576 18944 250626 19000
rect 250576 18942 250668 18944
rect 250621 18940 250668 18942
rect 250732 18940 250738 19004
rect 418654 18940 418660 19004
rect 418724 19002 418730 19004
rect 513414 19002 513420 19004
rect 418724 18942 513420 19002
rect 418724 18940 418730 18942
rect 513414 18940 513420 18942
rect 513484 18940 513490 19004
rect 515765 19002 515812 19004
rect 515720 19000 515812 19002
rect 515720 18944 515770 19000
rect 515720 18942 515812 18944
rect 515765 18940 515812 18942
rect 515876 18940 515882 19004
rect 247493 18939 247559 18940
rect 250621 18939 250687 18940
rect 515765 18939 515831 18940
rect 56041 18868 56107 18869
rect 55990 18804 55996 18868
rect 56060 18866 56107 18868
rect 58157 18868 58223 18869
rect 73705 18868 73771 18869
rect 58157 18866 58204 18868
rect 56060 18864 56152 18866
rect 56102 18808 56152 18864
rect 56060 18806 56152 18808
rect 58112 18864 58204 18866
rect 58112 18808 58162 18864
rect 58112 18806 58204 18808
rect 56060 18804 56107 18806
rect 56041 18803 56107 18804
rect 58157 18804 58204 18806
rect 58268 18804 58274 18868
rect 73654 18804 73660 18868
rect 73724 18866 73771 18868
rect 185485 18866 185551 18869
rect 252277 18868 252343 18869
rect 253565 18868 253631 18869
rect 238150 18866 238156 18868
rect 73724 18864 73816 18866
rect 73766 18808 73816 18864
rect 73724 18806 73816 18808
rect 185485 18864 238156 18866
rect 185485 18808 185490 18864
rect 185546 18808 238156 18864
rect 185485 18806 238156 18808
rect 73724 18804 73771 18806
rect 58157 18803 58223 18804
rect 73705 18803 73771 18804
rect 185485 18803 185551 18806
rect 238150 18804 238156 18806
rect 238220 18804 238226 18868
rect 252277 18866 252324 18868
rect 252232 18864 252324 18866
rect 252232 18808 252282 18864
rect 252232 18806 252324 18808
rect 252277 18804 252324 18806
rect 252388 18804 252394 18868
rect 253565 18866 253612 18868
rect 253520 18864 253612 18866
rect 253520 18808 253570 18864
rect 253520 18806 253612 18808
rect 253565 18804 253612 18806
rect 253676 18804 253682 18868
rect 399661 18866 399727 18869
rect 470869 18868 470935 18869
rect 465942 18866 465948 18868
rect 399661 18864 465948 18866
rect 399661 18808 399666 18864
rect 399722 18808 465948 18864
rect 399661 18806 465948 18808
rect 252277 18803 252343 18804
rect 253565 18803 253631 18804
rect 399661 18803 399727 18806
rect 465942 18804 465948 18806
rect 466012 18804 466018 18868
rect 470869 18866 470916 18868
rect 470824 18864 470916 18866
rect 470824 18808 470874 18864
rect 470824 18806 470916 18808
rect 470869 18804 470916 18806
rect 470980 18804 470986 18868
rect 485037 18866 485103 18869
rect 501045 18866 501111 18869
rect 505829 18868 505895 18869
rect 508405 18868 508471 18869
rect 505829 18866 505876 18868
rect 485037 18864 501111 18866
rect 485037 18808 485042 18864
rect 485098 18808 501050 18864
rect 501106 18808 501111 18864
rect 485037 18806 501111 18808
rect 505784 18864 505876 18866
rect 505784 18808 505834 18864
rect 505784 18806 505876 18808
rect 470869 18803 470935 18804
rect 485037 18803 485103 18806
rect 501045 18803 501111 18806
rect 505829 18804 505876 18806
rect 505940 18804 505946 18868
rect 508405 18866 508452 18868
rect 508360 18864 508452 18866
rect 508360 18808 508410 18864
rect 508360 18806 508452 18808
rect 508405 18804 508452 18806
rect 508516 18804 508522 18868
rect 505829 18803 505895 18804
rect 508405 18803 508471 18804
rect 50889 18732 50955 18733
rect 53649 18732 53715 18733
rect 50838 18668 50844 18732
rect 50908 18730 50955 18732
rect 50908 18728 51000 18730
rect 50950 18672 51000 18728
rect 50908 18670 51000 18672
rect 50908 18668 50955 18670
rect 53598 18668 53604 18732
rect 53668 18730 53715 18732
rect 188889 18730 188955 18733
rect 255957 18732 256023 18733
rect 258349 18732 258415 18733
rect 237046 18730 237052 18732
rect 53668 18728 53760 18730
rect 53710 18672 53760 18728
rect 53668 18670 53760 18672
rect 188889 18728 237052 18730
rect 188889 18672 188894 18728
rect 188950 18672 237052 18728
rect 188889 18670 237052 18672
rect 53668 18668 53715 18670
rect 50889 18667 50955 18668
rect 53649 18667 53715 18668
rect 188889 18667 188955 18670
rect 237046 18668 237052 18670
rect 237116 18668 237122 18732
rect 255957 18730 256004 18732
rect 255912 18728 256004 18730
rect 255912 18672 255962 18728
rect 255912 18670 256004 18672
rect 255957 18668 256004 18670
rect 256068 18668 256074 18732
rect 258349 18730 258396 18732
rect 258304 18728 258396 18730
rect 258304 18672 258354 18728
rect 258304 18670 258396 18672
rect 258349 18668 258396 18670
rect 258460 18668 258466 18732
rect 402237 18730 402303 18733
rect 523309 18732 523375 18733
rect 525885 18732 525951 18733
rect 523309 18730 523356 18732
rect 402237 18728 451290 18730
rect 402237 18672 402242 18728
rect 402298 18672 451290 18728
rect 402237 18670 451290 18672
rect 523264 18728 523356 18730
rect 523264 18672 523314 18728
rect 523264 18670 523356 18672
rect 255957 18667 256023 18668
rect 258349 18667 258415 18668
rect 402237 18667 402303 18670
rect 106089 18596 106155 18597
rect 108665 18596 108731 18597
rect 235993 18596 236059 18597
rect 106038 18532 106044 18596
rect 106108 18594 106155 18596
rect 106108 18592 106200 18594
rect 106150 18536 106200 18592
rect 106108 18534 106200 18536
rect 106108 18532 106155 18534
rect 108614 18532 108620 18596
rect 108684 18594 108731 18596
rect 108684 18592 108776 18594
rect 108726 18536 108776 18592
rect 108684 18534 108776 18536
rect 108684 18532 108731 18534
rect 235942 18532 235948 18596
rect 236012 18594 236059 18596
rect 243077 18596 243143 18597
rect 243077 18594 243124 18596
rect 236012 18592 236104 18594
rect 236054 18536 236104 18592
rect 236012 18534 236104 18536
rect 243032 18592 243124 18594
rect 243032 18536 243082 18592
rect 243032 18534 243124 18536
rect 236012 18532 236059 18534
rect 106089 18531 106155 18532
rect 108665 18531 108731 18532
rect 235993 18531 236059 18532
rect 243077 18532 243124 18534
rect 243188 18532 243194 18596
rect 451230 18594 451290 18670
rect 523309 18668 523356 18670
rect 523420 18668 523426 18732
rect 525885 18730 525932 18732
rect 525840 18728 525932 18730
rect 525840 18672 525890 18728
rect 525840 18670 525932 18672
rect 525885 18668 525932 18670
rect 525996 18668 526002 18732
rect 523309 18667 523375 18668
rect 525885 18667 525951 18668
rect 463550 18594 463556 18596
rect 451230 18534 463556 18594
rect 463550 18532 463556 18534
rect 463620 18532 463626 18596
rect 243077 18531 243143 18532
rect 113449 18460 113515 18461
rect 113398 18396 113404 18460
rect 113468 18458 113515 18460
rect 113468 18456 113560 18458
rect 113510 18400 113560 18456
rect 113468 18398 113560 18400
rect 113468 18396 113515 18398
rect 113449 18395 113515 18396
rect 41638 18124 41644 18188
rect 41708 18124 41714 18188
rect 45318 18124 45324 18188
rect 45388 18124 45394 18188
rect 74390 18124 74396 18188
rect 74460 18124 74466 18188
rect 36537 17914 36603 17917
rect 37038 17914 37044 17916
rect 36537 17912 37044 17914
rect 36537 17856 36542 17912
rect 36598 17856 37044 17912
rect 36537 17854 37044 17856
rect 36537 17851 36603 17854
rect 37038 17852 37044 17854
rect 37108 17852 37114 17916
rect 19006 17716 19012 17780
rect 19076 17778 19082 17780
rect 41646 17778 41706 18124
rect 45326 17917 45386 18124
rect 43069 17916 43135 17917
rect 44173 17916 44239 17917
rect 43069 17912 43116 17916
rect 43180 17914 43186 17916
rect 43069 17856 43074 17912
rect 43069 17852 43116 17856
rect 43180 17854 43226 17914
rect 44173 17912 44220 17916
rect 44284 17914 44290 17916
rect 44173 17856 44178 17912
rect 43180 17852 43186 17854
rect 44173 17852 44220 17856
rect 44284 17854 44330 17914
rect 45326 17912 45435 17917
rect 46657 17916 46723 17917
rect 47577 17916 47643 17917
rect 48681 17916 48747 17917
rect 50153 17916 50219 17917
rect 51441 17916 51507 17917
rect 59537 17916 59603 17917
rect 46606 17914 46612 17916
rect 45326 17856 45374 17912
rect 45430 17856 45435 17912
rect 45326 17854 45435 17856
rect 46566 17854 46612 17914
rect 46676 17912 46723 17916
rect 47526 17914 47532 17916
rect 46718 17856 46723 17912
rect 44284 17852 44290 17854
rect 43069 17851 43135 17852
rect 44173 17851 44239 17852
rect 45369 17851 45435 17854
rect 46606 17852 46612 17854
rect 46676 17852 46723 17856
rect 47486 17854 47532 17914
rect 47596 17912 47643 17916
rect 48630 17914 48636 17916
rect 47638 17856 47643 17912
rect 47526 17852 47532 17854
rect 47596 17852 47643 17856
rect 48590 17854 48636 17914
rect 48700 17912 48747 17916
rect 50102 17914 50108 17916
rect 48742 17856 48747 17912
rect 48630 17852 48636 17854
rect 48700 17852 48747 17856
rect 50062 17854 50108 17914
rect 50172 17912 50219 17916
rect 51390 17914 51396 17916
rect 50214 17856 50219 17912
rect 50102 17852 50108 17854
rect 50172 17852 50219 17856
rect 51350 17854 51396 17914
rect 51460 17912 51507 17916
rect 59486 17914 59492 17916
rect 51502 17856 51507 17912
rect 51390 17852 51396 17854
rect 51460 17852 51507 17856
rect 59446 17854 59492 17914
rect 59556 17912 59603 17916
rect 59598 17856 59603 17912
rect 59486 17852 59492 17854
rect 59556 17852 59603 17856
rect 46657 17851 46723 17852
rect 47577 17851 47643 17852
rect 48681 17851 48747 17852
rect 50153 17851 50219 17852
rect 51441 17851 51507 17852
rect 59537 17851 59603 17852
rect 60457 17914 60523 17917
rect 60590 17914 60596 17916
rect 60457 17912 60596 17914
rect 60457 17856 60462 17912
rect 60518 17856 60596 17912
rect 60457 17854 60596 17856
rect 60457 17851 60523 17854
rect 60590 17852 60596 17854
rect 60660 17852 60666 17916
rect 61142 17852 61148 17916
rect 61212 17914 61218 17916
rect 62021 17914 62087 17917
rect 61212 17912 62087 17914
rect 61212 17856 62026 17912
rect 62082 17856 62087 17912
rect 61212 17854 62087 17856
rect 61212 17852 61218 17854
rect 62021 17851 62087 17854
rect 63534 17852 63540 17916
rect 63604 17914 63610 17916
rect 64689 17914 64755 17917
rect 63604 17912 64755 17914
rect 63604 17856 64694 17912
rect 64750 17856 64755 17912
rect 63604 17854 64755 17856
rect 63604 17852 63610 17854
rect 64689 17851 64755 17854
rect 65926 17852 65932 17916
rect 65996 17914 66002 17916
rect 66161 17914 66227 17917
rect 65996 17912 66227 17914
rect 65996 17856 66166 17912
rect 66222 17856 66227 17912
rect 65996 17854 66227 17856
rect 65996 17852 66002 17854
rect 66161 17851 66227 17854
rect 67633 17914 67699 17917
rect 68686 17914 68692 17916
rect 67633 17912 68692 17914
rect 67633 17856 67638 17912
rect 67694 17856 68692 17912
rect 67633 17854 68692 17856
rect 67633 17851 67699 17854
rect 68686 17852 68692 17854
rect 68756 17852 68762 17916
rect 71773 17914 71839 17917
rect 72182 17914 72188 17916
rect 71773 17912 72188 17914
rect 71773 17856 71778 17912
rect 71834 17856 72188 17912
rect 71773 17854 72188 17856
rect 71773 17851 71839 17854
rect 72182 17852 72188 17854
rect 72252 17852 72258 17916
rect 73153 17914 73219 17917
rect 74398 17914 74458 18124
rect 458357 18052 458423 18053
rect 458357 18050 458404 18052
rect 458312 18048 458404 18050
rect 458312 17992 458362 18048
rect 458312 17990 458404 17992
rect 458357 17988 458404 17990
rect 458468 17988 458474 18052
rect 458357 17987 458423 17988
rect 73153 17912 74458 17914
rect 73153 17856 73158 17912
rect 73214 17856 74458 17912
rect 73153 17854 74458 17856
rect 73153 17851 73219 17854
rect 78438 17852 78444 17916
rect 78508 17914 78514 17916
rect 78581 17914 78647 17917
rect 125961 17916 126027 17917
rect 78508 17912 78647 17914
rect 78508 17856 78586 17912
rect 78642 17856 78647 17912
rect 78508 17854 78647 17856
rect 78508 17852 78514 17854
rect 78581 17851 78647 17854
rect 125910 17852 125916 17916
rect 125980 17914 126027 17916
rect 268326 17914 268332 17916
rect 125980 17912 126072 17914
rect 126022 17856 126072 17912
rect 125980 17854 126072 17856
rect 258030 17854 268332 17914
rect 125980 17852 126027 17854
rect 125961 17851 126027 17852
rect 19076 17718 41706 17778
rect 19076 17716 19082 17718
rect 48262 17716 48268 17780
rect 48332 17778 48338 17780
rect 181437 17778 181503 17781
rect 48332 17776 181503 17778
rect 48332 17720 181442 17776
rect 181498 17720 181503 17776
rect 48332 17718 181503 17720
rect 48332 17716 48338 17718
rect 181437 17715 181503 17718
rect 192334 17716 192340 17780
rect 192404 17778 192410 17780
rect 258030 17778 258090 17854
rect 268326 17852 268332 17854
rect 268396 17852 268402 17916
rect 273253 17914 273319 17917
rect 273478 17914 273484 17916
rect 273253 17912 273484 17914
rect 273253 17856 273258 17912
rect 273314 17856 273484 17912
rect 273253 17854 273484 17856
rect 273253 17851 273319 17854
rect 273478 17852 273484 17854
rect 273548 17852 273554 17916
rect 277158 17852 277164 17916
rect 277228 17914 277234 17916
rect 277393 17914 277459 17917
rect 277228 17912 277459 17914
rect 277228 17856 277398 17912
rect 277454 17856 277459 17912
rect 277228 17854 277459 17856
rect 277228 17852 277234 17854
rect 277393 17851 277459 17854
rect 280153 17914 280219 17917
rect 436093 17916 436159 17917
rect 280838 17914 280844 17916
rect 280153 17912 280844 17914
rect 280153 17856 280158 17912
rect 280214 17856 280844 17912
rect 280153 17854 280844 17856
rect 280153 17851 280219 17854
rect 280838 17852 280844 17854
rect 280908 17852 280914 17916
rect 436093 17914 436140 17916
rect 436048 17912 436140 17914
rect 436048 17856 436098 17912
rect 436048 17854 436140 17856
rect 436093 17852 436140 17854
rect 436204 17852 436210 17916
rect 436277 17914 436343 17917
rect 437054 17914 437060 17916
rect 436277 17912 437060 17914
rect 436277 17856 436282 17912
rect 436338 17856 437060 17912
rect 436277 17854 437060 17856
rect 436093 17851 436159 17852
rect 436277 17851 436343 17854
rect 437054 17852 437060 17854
rect 437124 17852 437130 17916
rect 437473 17914 437539 17917
rect 438342 17914 438348 17916
rect 437473 17912 438348 17914
rect 437473 17856 437478 17912
rect 437534 17856 438348 17912
rect 437473 17854 438348 17856
rect 437473 17851 437539 17854
rect 438342 17852 438348 17854
rect 438412 17852 438418 17916
rect 438853 17914 438919 17917
rect 439630 17914 439636 17916
rect 438853 17912 439636 17914
rect 438853 17856 438858 17912
rect 438914 17856 439636 17912
rect 438853 17854 439636 17856
rect 438853 17851 438919 17854
rect 439630 17852 439636 17854
rect 439700 17852 439706 17916
rect 440233 17914 440299 17917
rect 440550 17914 440556 17916
rect 440233 17912 440556 17914
rect 440233 17856 440238 17912
rect 440294 17856 440556 17912
rect 440233 17854 440556 17856
rect 440233 17851 440299 17854
rect 440550 17852 440556 17854
rect 440620 17852 440626 17916
rect 441705 17914 441771 17917
rect 443085 17916 443151 17917
rect 444281 17916 444347 17917
rect 442022 17914 442028 17916
rect 441705 17912 442028 17914
rect 441705 17856 441710 17912
rect 441766 17856 442028 17912
rect 441705 17854 442028 17856
rect 441705 17851 441771 17854
rect 442022 17852 442028 17854
rect 442092 17852 442098 17916
rect 443085 17912 443132 17916
rect 443196 17914 443202 17916
rect 444230 17914 444236 17916
rect 443085 17856 443090 17912
rect 443085 17852 443132 17856
rect 443196 17854 443242 17914
rect 444190 17854 444236 17914
rect 444300 17912 444347 17916
rect 444342 17856 444347 17912
rect 443196 17852 443202 17854
rect 444230 17852 444236 17854
rect 444300 17852 444347 17856
rect 443085 17851 443151 17852
rect 444281 17851 444347 17852
rect 445661 17916 445727 17917
rect 446489 17916 446555 17917
rect 445661 17912 445708 17916
rect 445772 17914 445778 17916
rect 446438 17914 446444 17916
rect 445661 17856 445666 17912
rect 445661 17852 445708 17856
rect 445772 17854 445818 17914
rect 446398 17854 446444 17914
rect 446508 17912 446555 17916
rect 446550 17856 446555 17912
rect 445772 17852 445778 17854
rect 446438 17852 446444 17854
rect 446508 17852 446555 17856
rect 445661 17851 445727 17852
rect 446489 17851 446555 17852
rect 447133 17914 447199 17917
rect 448278 17914 448284 17916
rect 447133 17912 448284 17914
rect 447133 17856 447138 17912
rect 447194 17856 448284 17912
rect 447133 17854 448284 17856
rect 447133 17851 447199 17854
rect 448278 17852 448284 17854
rect 448348 17852 448354 17916
rect 449893 17914 449959 17917
rect 450670 17914 450676 17916
rect 449893 17912 450676 17914
rect 449893 17856 449898 17912
rect 449954 17856 450676 17912
rect 449893 17854 450676 17856
rect 449893 17851 449959 17854
rect 450670 17852 450676 17854
rect 450740 17852 450746 17916
rect 451273 17914 451339 17917
rect 452285 17916 452351 17917
rect 453481 17916 453547 17917
rect 451406 17914 451412 17916
rect 451273 17912 451412 17914
rect 451273 17856 451278 17912
rect 451334 17856 451412 17912
rect 451273 17854 451412 17856
rect 451273 17851 451339 17854
rect 451406 17852 451412 17854
rect 451476 17852 451482 17916
rect 452285 17912 452332 17916
rect 452396 17914 452402 17916
rect 453430 17914 453436 17916
rect 452285 17856 452290 17912
rect 452285 17852 452332 17856
rect 452396 17854 452442 17914
rect 453390 17854 453436 17914
rect 453500 17912 453547 17916
rect 453542 17856 453547 17912
rect 452396 17852 452402 17854
rect 453430 17852 453436 17854
rect 453500 17852 453547 17856
rect 452285 17851 452351 17852
rect 453481 17851 453547 17852
rect 454033 17914 454099 17917
rect 454534 17914 454540 17916
rect 454033 17912 454540 17914
rect 454033 17856 454038 17912
rect 454094 17856 454540 17912
rect 454033 17854 454540 17856
rect 454033 17851 454099 17854
rect 454534 17852 454540 17854
rect 454604 17852 454610 17916
rect 455413 17914 455479 17917
rect 456006 17914 456012 17916
rect 455413 17912 456012 17914
rect 455413 17856 455418 17912
rect 455474 17856 456012 17912
rect 455413 17854 456012 17856
rect 455413 17851 455479 17854
rect 456006 17852 456012 17854
rect 456076 17852 456082 17916
rect 457110 17852 457116 17916
rect 457180 17914 457186 17916
rect 457345 17914 457411 17917
rect 458081 17916 458147 17917
rect 458030 17914 458036 17916
rect 457180 17912 457411 17914
rect 457180 17856 457350 17912
rect 457406 17856 457411 17912
rect 457180 17854 457411 17856
rect 457990 17854 458036 17914
rect 458100 17912 458147 17916
rect 458142 17856 458147 17912
rect 457180 17852 457186 17854
rect 457345 17851 457411 17854
rect 458030 17852 458036 17854
rect 458100 17852 458147 17856
rect 458081 17851 458147 17852
rect 458265 17914 458331 17917
rect 459318 17914 459324 17916
rect 458265 17912 459324 17914
rect 458265 17856 458270 17912
rect 458326 17856 459324 17912
rect 458265 17854 459324 17856
rect 458265 17851 458331 17854
rect 459318 17852 459324 17854
rect 459388 17852 459394 17916
rect 459461 17914 459527 17917
rect 461710 17914 461716 17916
rect 459461 17912 461716 17914
rect 459461 17856 459466 17912
rect 459522 17856 461716 17912
rect 459461 17854 461716 17856
rect 459461 17851 459527 17854
rect 461710 17852 461716 17854
rect 461780 17852 461786 17916
rect 462313 17914 462379 17917
rect 462814 17914 462820 17916
rect 462313 17912 462820 17914
rect 462313 17856 462318 17912
rect 462374 17856 462820 17912
rect 462313 17854 462820 17856
rect 462313 17851 462379 17854
rect 462814 17852 462820 17854
rect 462884 17852 462890 17916
rect 463693 17914 463759 17917
rect 463918 17914 463924 17916
rect 463693 17912 463924 17914
rect 463693 17856 463698 17912
rect 463754 17856 463924 17912
rect 463693 17854 463924 17856
rect 463693 17851 463759 17854
rect 463918 17852 463924 17854
rect 463988 17852 463994 17916
rect 465073 17914 465139 17917
rect 466310 17914 466316 17916
rect 465073 17912 466316 17914
rect 465073 17856 465078 17912
rect 465134 17856 466316 17912
rect 465073 17854 466316 17856
rect 465073 17851 465139 17854
rect 466310 17852 466316 17854
rect 466380 17852 466386 17916
rect 466453 17914 466519 17917
rect 467598 17914 467604 17916
rect 466453 17912 467604 17914
rect 466453 17856 466458 17912
rect 466514 17856 467604 17912
rect 466453 17854 467604 17856
rect 466453 17851 466519 17854
rect 467598 17852 467604 17854
rect 467668 17852 467674 17916
rect 467833 17914 467899 17917
rect 468702 17914 468708 17916
rect 467833 17912 468708 17914
rect 467833 17856 467838 17912
rect 467894 17856 468708 17912
rect 467833 17854 468708 17856
rect 467833 17851 467899 17854
rect 468702 17852 468708 17854
rect 468772 17852 468778 17916
rect 473353 17914 473419 17917
rect 474406 17914 474412 17916
rect 473353 17912 474412 17914
rect 473353 17856 473358 17912
rect 473414 17856 474412 17912
rect 473353 17854 474412 17856
rect 473353 17851 473419 17854
rect 474406 17852 474412 17854
rect 474476 17852 474482 17916
rect 476113 17914 476179 17917
rect 476982 17914 476988 17916
rect 476113 17912 476988 17914
rect 476113 17856 476118 17912
rect 476174 17856 476988 17912
rect 476113 17854 476988 17856
rect 476113 17851 476179 17854
rect 476982 17852 476988 17854
rect 477052 17852 477058 17916
rect 478873 17914 478939 17917
rect 479190 17914 479196 17916
rect 478873 17912 479196 17914
rect 478873 17856 478878 17912
rect 478934 17856 479196 17912
rect 478873 17854 479196 17856
rect 478873 17851 478939 17854
rect 479190 17852 479196 17854
rect 479260 17852 479266 17916
rect 263593 17780 263659 17781
rect 192404 17718 258090 17778
rect 192404 17716 192410 17718
rect 263542 17716 263548 17780
rect 263612 17778 263659 17780
rect 264973 17778 265039 17781
rect 265934 17778 265940 17780
rect 263612 17776 263704 17778
rect 263654 17720 263704 17776
rect 263612 17718 263704 17720
rect 264973 17776 265940 17778
rect 264973 17720 264978 17776
rect 265034 17720 265940 17776
rect 264973 17718 265940 17720
rect 263612 17716 263659 17718
rect 263593 17715 263659 17716
rect 264973 17715 265039 17718
rect 265934 17716 265940 17718
rect 266004 17716 266010 17780
rect 388437 17778 388503 17781
rect 473302 17778 473308 17780
rect 388437 17776 473308 17778
rect 388437 17720 388442 17776
rect 388498 17720 473308 17776
rect 388437 17718 473308 17720
rect 388437 17715 388503 17718
rect 473302 17716 473308 17718
rect 473372 17716 473378 17780
rect 475377 17778 475443 17781
rect 480662 17778 480668 17780
rect 475377 17776 480668 17778
rect 475377 17720 475382 17776
rect 475438 17720 480668 17776
rect 475377 17718 480668 17720
rect 475377 17715 475443 17718
rect 480662 17716 480668 17718
rect 480732 17716 480738 17780
rect 19793 17642 19859 17645
rect 40534 17642 40540 17644
rect 19793 17640 40540 17642
rect 19793 17584 19798 17640
rect 19854 17584 40540 17640
rect 19793 17582 40540 17584
rect 19793 17579 19859 17582
rect 40534 17580 40540 17582
rect 40604 17580 40610 17644
rect 53833 17642 53899 17645
rect 54518 17642 54524 17644
rect 53833 17640 54524 17642
rect 53833 17584 53838 17640
rect 53894 17584 54524 17640
rect 53833 17582 54524 17584
rect 53833 17579 53899 17582
rect 54518 17580 54524 17582
rect 54588 17642 54594 17644
rect 68185 17642 68251 17645
rect 54588 17640 68251 17642
rect 54588 17584 68190 17640
rect 68246 17584 68251 17640
rect 54588 17582 68251 17584
rect 54588 17580 54594 17582
rect 68185 17579 68251 17582
rect 68318 17580 68324 17644
rect 68388 17642 68394 17644
rect 68921 17642 68987 17645
rect 68388 17640 68987 17642
rect 68388 17584 68926 17640
rect 68982 17584 68987 17640
rect 68388 17582 68987 17584
rect 68388 17580 68394 17582
rect 68921 17579 68987 17582
rect 70393 17642 70459 17645
rect 71262 17642 71268 17644
rect 70393 17640 71268 17642
rect 70393 17584 70398 17640
rect 70454 17584 71268 17640
rect 70393 17582 71268 17584
rect 70393 17579 70459 17582
rect 71262 17580 71268 17582
rect 71332 17580 71338 17644
rect 83590 17580 83596 17644
rect 83660 17642 83666 17644
rect 83825 17642 83891 17645
rect 83660 17640 83891 17642
rect 83660 17584 83830 17640
rect 83886 17584 83891 17640
rect 83660 17582 83891 17584
rect 83660 17580 83666 17582
rect 83825 17579 83891 17582
rect 115790 17580 115796 17644
rect 115860 17642 115866 17644
rect 188286 17642 188292 17644
rect 115860 17582 188292 17642
rect 115860 17580 115866 17582
rect 188286 17580 188292 17582
rect 188356 17580 188362 17644
rect 192518 17580 192524 17644
rect 192588 17642 192594 17644
rect 254526 17642 254532 17644
rect 192588 17582 254532 17642
rect 192588 17580 192594 17582
rect 254526 17580 254532 17582
rect 254596 17580 254602 17644
rect 259545 17642 259611 17645
rect 260598 17642 260604 17644
rect 259545 17640 260604 17642
rect 259545 17584 259550 17640
rect 259606 17584 260604 17640
rect 259545 17582 260604 17584
rect 259545 17579 259611 17582
rect 260598 17580 260604 17582
rect 260668 17580 260674 17644
rect 260833 17642 260899 17645
rect 260966 17642 260972 17644
rect 260833 17640 260972 17642
rect 260833 17584 260838 17640
rect 260894 17584 260972 17640
rect 260833 17582 260972 17584
rect 260833 17579 260899 17582
rect 260966 17580 260972 17582
rect 261036 17580 261042 17644
rect 270493 17642 270559 17645
rect 270902 17642 270908 17644
rect 270493 17640 270908 17642
rect 270493 17584 270498 17640
rect 270554 17584 270908 17640
rect 270493 17582 270908 17584
rect 270493 17579 270559 17582
rect 270902 17580 270908 17582
rect 270972 17580 270978 17644
rect 404997 17642 405063 17645
rect 483422 17642 483428 17644
rect 404997 17640 483428 17642
rect 404997 17584 405002 17640
rect 405058 17584 483428 17640
rect 404997 17582 483428 17584
rect 404997 17579 405063 17582
rect 483422 17580 483428 17582
rect 483492 17580 483498 17644
rect 19149 17506 19215 17509
rect 38510 17506 38516 17508
rect 19149 17504 38516 17506
rect 19149 17448 19154 17504
rect 19210 17448 38516 17504
rect 19149 17446 38516 17448
rect 19149 17443 19215 17446
rect 38510 17444 38516 17446
rect 38580 17444 38586 17508
rect 58198 17444 58204 17508
rect 58268 17506 58274 17508
rect 69657 17506 69723 17509
rect 58268 17504 69723 17506
rect 58268 17448 69662 17504
rect 69718 17448 69723 17504
rect 58268 17446 69723 17448
rect 58268 17444 58274 17446
rect 69657 17443 69723 17446
rect 75913 17506 75979 17509
rect 76966 17506 76972 17508
rect 75913 17504 76972 17506
rect 75913 17448 75918 17504
rect 75974 17448 76972 17504
rect 75913 17446 76972 17448
rect 75913 17443 75979 17446
rect 76966 17444 76972 17446
rect 77036 17444 77042 17508
rect 78673 17506 78739 17509
rect 88241 17508 88307 17509
rect 93577 17508 93643 17509
rect 79174 17506 79180 17508
rect 78673 17504 79180 17506
rect 78673 17448 78678 17504
rect 78734 17448 79180 17504
rect 78673 17446 79180 17448
rect 78673 17443 78739 17446
rect 79174 17444 79180 17446
rect 79244 17444 79250 17508
rect 88190 17444 88196 17508
rect 88260 17506 88307 17508
rect 88260 17504 88352 17506
rect 88302 17448 88352 17504
rect 88260 17446 88352 17448
rect 88260 17444 88307 17446
rect 93526 17444 93532 17508
rect 93596 17506 93643 17508
rect 93596 17504 93688 17506
rect 93638 17448 93688 17504
rect 93596 17446 93688 17448
rect 93596 17444 93643 17446
rect 122598 17444 122604 17508
rect 122668 17506 122674 17508
rect 191046 17506 191052 17508
rect 122668 17446 191052 17506
rect 122668 17444 122674 17446
rect 191046 17444 191052 17446
rect 191116 17444 191122 17508
rect 191373 17506 191439 17509
rect 259453 17508 259519 17509
rect 253422 17506 253428 17508
rect 191373 17504 253428 17506
rect 191373 17448 191378 17504
rect 191434 17448 253428 17504
rect 191373 17446 253428 17448
rect 88241 17443 88307 17444
rect 93577 17443 93643 17444
rect 191373 17443 191439 17446
rect 253422 17444 253428 17446
rect 253492 17444 253498 17508
rect 259453 17506 259500 17508
rect 259408 17504 259500 17506
rect 259408 17448 259458 17504
rect 259408 17446 259500 17448
rect 259453 17444 259500 17446
rect 259564 17444 259570 17508
rect 405181 17506 405247 17509
rect 475377 17506 475443 17509
rect 405181 17504 475443 17506
rect 405181 17448 405186 17504
rect 405242 17448 475382 17504
rect 475438 17448 475443 17504
rect 405181 17446 475443 17448
rect 259453 17443 259519 17444
rect 405181 17443 405247 17446
rect 475377 17443 475443 17446
rect 18689 17370 18755 17373
rect 56910 17370 56916 17372
rect 18689 17368 56916 17370
rect 18689 17312 18694 17368
rect 18750 17312 56916 17368
rect 18689 17310 56916 17312
rect 18689 17307 18755 17310
rect 56910 17308 56916 17310
rect 56980 17370 56986 17372
rect 57881 17370 57947 17373
rect 56980 17368 57947 17370
rect 56980 17312 57886 17368
rect 57942 17312 57947 17368
rect 56980 17310 57947 17312
rect 56980 17308 56986 17310
rect 57881 17307 57947 17310
rect 65057 17370 65123 17373
rect 66253 17372 66319 17373
rect 67633 17372 67699 17373
rect 65190 17370 65196 17372
rect 65057 17368 65196 17370
rect 65057 17312 65062 17368
rect 65118 17312 65196 17368
rect 65057 17310 65196 17312
rect 65057 17307 65123 17310
rect 65190 17308 65196 17310
rect 65260 17308 65266 17372
rect 66253 17370 66300 17372
rect 66208 17368 66300 17370
rect 66208 17312 66258 17368
rect 66208 17310 66300 17312
rect 66253 17308 66300 17310
rect 66364 17308 66370 17372
rect 67582 17308 67588 17372
rect 67652 17370 67699 17372
rect 68185 17370 68251 17373
rect 73286 17370 73292 17372
rect 67652 17368 67744 17370
rect 67694 17312 67744 17368
rect 67652 17310 67744 17312
rect 68185 17368 73292 17370
rect 68185 17312 68190 17368
rect 68246 17312 73292 17368
rect 68185 17310 73292 17312
rect 67652 17308 67699 17310
rect 66253 17307 66319 17308
rect 67633 17307 67699 17308
rect 68185 17307 68251 17310
rect 73286 17308 73292 17310
rect 73356 17308 73362 17372
rect 98494 17308 98500 17372
rect 98564 17370 98570 17372
rect 99281 17370 99347 17373
rect 98564 17368 99347 17370
rect 98564 17312 99286 17368
rect 99342 17312 99347 17368
rect 98564 17310 99347 17312
rect 98564 17308 98570 17310
rect 99281 17307 99347 17310
rect 111006 17308 111012 17372
rect 111076 17370 111082 17372
rect 111701 17370 111767 17373
rect 111076 17368 111767 17370
rect 111076 17312 111706 17368
rect 111762 17312 111767 17368
rect 111076 17310 111767 17312
rect 111076 17308 111082 17310
rect 111701 17307 111767 17310
rect 187417 17370 187483 17373
rect 248638 17370 248644 17372
rect 187417 17368 248644 17370
rect 187417 17312 187422 17368
rect 187478 17312 248644 17368
rect 187417 17310 248644 17312
rect 187417 17307 187483 17310
rect 248638 17308 248644 17310
rect 248708 17308 248714 17372
rect 255313 17370 255379 17373
rect 255814 17370 255820 17372
rect 255313 17368 255820 17370
rect 255313 17312 255318 17368
rect 255374 17312 255820 17368
rect 255313 17310 255820 17312
rect 255313 17307 255379 17310
rect 255814 17308 255820 17310
rect 255884 17308 255890 17372
rect 256693 17370 256759 17373
rect 256918 17370 256924 17372
rect 256693 17368 256924 17370
rect 256693 17312 256698 17368
rect 256754 17312 256924 17368
rect 256693 17310 256924 17312
rect 256693 17307 256759 17310
rect 256918 17308 256924 17310
rect 256988 17308 256994 17372
rect 258073 17370 258139 17373
rect 258390 17370 258396 17372
rect 258073 17368 258396 17370
rect 258073 17312 258078 17368
rect 258134 17312 258396 17368
rect 258073 17310 258396 17312
rect 258073 17307 258139 17310
rect 258390 17308 258396 17310
rect 258460 17308 258466 17372
rect 407757 17370 407823 17373
rect 471697 17370 471763 17373
rect 476062 17370 476068 17372
rect 407757 17368 471763 17370
rect 407757 17312 407762 17368
rect 407818 17312 471702 17368
rect 471758 17312 471763 17368
rect 407757 17310 471763 17312
rect 407757 17307 407823 17310
rect 471697 17307 471763 17310
rect 471838 17310 476068 17370
rect 18965 17234 19031 17237
rect 35934 17234 35940 17236
rect 18965 17232 35940 17234
rect 18965 17176 18970 17232
rect 19026 17176 35940 17232
rect 18965 17174 35940 17176
rect 18965 17171 19031 17174
rect 35934 17172 35940 17174
rect 36004 17172 36010 17236
rect 38653 17234 38719 17237
rect 39614 17234 39620 17236
rect 38653 17232 39620 17234
rect 38653 17176 38658 17232
rect 38714 17176 39620 17232
rect 38653 17174 39620 17176
rect 38653 17171 38719 17174
rect 39614 17172 39620 17174
rect 39684 17172 39690 17236
rect 60733 17234 60799 17237
rect 61694 17234 61700 17236
rect 60733 17232 61700 17234
rect 60733 17176 60738 17232
rect 60794 17176 61700 17232
rect 60733 17174 61700 17176
rect 60733 17171 60799 17174
rect 61694 17172 61700 17174
rect 61764 17172 61770 17236
rect 62113 17234 62179 17237
rect 62798 17234 62804 17236
rect 62113 17232 62804 17234
rect 62113 17176 62118 17232
rect 62174 17176 62804 17232
rect 62113 17174 62804 17176
rect 62113 17171 62179 17174
rect 62798 17172 62804 17174
rect 62868 17172 62874 17236
rect 63493 17234 63559 17237
rect 63902 17234 63908 17236
rect 63493 17232 63908 17234
rect 63493 17176 63498 17232
rect 63554 17176 63908 17232
rect 63493 17174 63908 17176
rect 63493 17171 63559 17174
rect 63902 17172 63908 17174
rect 63972 17172 63978 17236
rect 69013 17234 69079 17237
rect 69790 17234 69796 17236
rect 69013 17232 69796 17234
rect 69013 17176 69018 17232
rect 69074 17176 69796 17232
rect 69013 17174 69796 17176
rect 69013 17171 69079 17174
rect 69790 17172 69796 17174
rect 69860 17172 69866 17236
rect 70894 17172 70900 17236
rect 70964 17234 70970 17236
rect 71681 17234 71747 17237
rect 70964 17232 71747 17234
rect 70964 17176 71686 17232
rect 71742 17176 71747 17232
rect 70964 17174 71747 17176
rect 70964 17172 70970 17174
rect 71681 17171 71747 17174
rect 74809 17234 74875 17237
rect 75678 17234 75684 17236
rect 74809 17232 75684 17234
rect 74809 17176 74814 17232
rect 74870 17176 75684 17232
rect 74809 17174 75684 17176
rect 74809 17171 74875 17174
rect 75678 17172 75684 17174
rect 75748 17172 75754 17236
rect 192702 17172 192708 17236
rect 192772 17234 192778 17236
rect 276054 17234 276060 17236
rect 192772 17174 276060 17234
rect 192772 17172 192778 17174
rect 276054 17172 276060 17174
rect 276124 17172 276130 17236
rect 282913 17234 282979 17237
rect 283414 17234 283420 17236
rect 282913 17232 283420 17234
rect 282913 17176 282918 17232
rect 282974 17176 283420 17232
rect 282913 17174 283420 17176
rect 282913 17171 282979 17174
rect 283414 17172 283420 17174
rect 283484 17172 283490 17236
rect 407941 17234 408007 17237
rect 471838 17234 471898 17310
rect 476062 17308 476068 17310
rect 476132 17308 476138 17372
rect 407941 17232 471898 17234
rect 407941 17176 407946 17232
rect 408002 17176 471898 17232
rect 407941 17174 471898 17176
rect 471973 17234 472039 17237
rect 472198 17234 472204 17236
rect 471973 17232 472204 17234
rect 471973 17176 471978 17232
rect 472034 17176 472204 17232
rect 471973 17174 472204 17176
rect 407941 17171 408007 17174
rect 471973 17171 472039 17174
rect 472198 17172 472204 17174
rect 472268 17172 472274 17236
rect 474733 17234 474799 17237
rect 475694 17234 475700 17236
rect 474733 17232 475700 17234
rect 474733 17176 474738 17232
rect 474794 17176 475700 17232
rect 474733 17174 475700 17176
rect 474733 17171 474799 17174
rect 475694 17172 475700 17174
rect 475764 17172 475770 17236
rect 251173 17100 251239 17101
rect 58566 17036 58572 17100
rect 58636 17098 58642 17100
rect 191782 17098 191788 17100
rect 58636 17038 191788 17098
rect 58636 17036 58642 17038
rect 191782 17036 191788 17038
rect 191852 17036 191858 17100
rect 251173 17098 251220 17100
rect 251128 17096 251220 17098
rect 251128 17040 251178 17096
rect 251128 17038 251220 17040
rect 251173 17036 251220 17038
rect 251284 17036 251290 17100
rect 414606 17036 414612 17100
rect 414676 17098 414682 17100
rect 465073 17098 465139 17101
rect 465206 17098 465212 17100
rect 414676 17038 431970 17098
rect 414676 17036 414682 17038
rect 251173 17035 251239 17036
rect 77293 16962 77359 16965
rect 78254 16962 78260 16964
rect 77293 16960 78260 16962
rect 77293 16904 77298 16960
rect 77354 16904 78260 16960
rect 77293 16902 78260 16904
rect 77293 16899 77359 16902
rect 78254 16900 78260 16902
rect 78324 16900 78330 16964
rect 431910 16962 431970 17038
rect 465073 17096 465212 17098
rect 465073 17040 465078 17096
rect 465134 17040 465212 17096
rect 465073 17038 465212 17040
rect 465073 17035 465139 17038
rect 465206 17036 465212 17038
rect 465276 17036 465282 17100
rect 469305 17098 469371 17101
rect 469622 17098 469628 17100
rect 469305 17096 469628 17098
rect 469305 17040 469310 17096
rect 469366 17040 469628 17096
rect 469305 17038 469628 17040
rect 469305 17035 469371 17038
rect 469622 17036 469628 17038
rect 469692 17036 469698 17100
rect 471697 17098 471763 17101
rect 478454 17098 478460 17100
rect 471697 17096 478460 17098
rect 471697 17040 471702 17096
rect 471758 17040 478460 17096
rect 471697 17038 478460 17040
rect 471697 17035 471763 17038
rect 478454 17036 478460 17038
rect 478524 17036 478530 17100
rect 453614 16962 453620 16964
rect 431910 16902 453620 16962
rect 453614 16900 453620 16902
rect 453684 16900 453690 16964
rect 477493 16962 477559 16965
rect 478086 16962 478092 16964
rect 477493 16960 478092 16962
rect 477493 16904 477498 16960
rect 477554 16904 478092 16960
rect 477493 16902 478092 16904
rect 477493 16899 477559 16902
rect 478086 16900 478092 16902
rect 478156 16900 478162 16964
rect 470869 16826 470935 16829
rect 471278 16826 471284 16828
rect 470869 16824 471284 16826
rect 470869 16768 470874 16824
rect 470930 16768 471284 16824
rect 470869 16766 471284 16768
rect 470869 16763 470935 16766
rect 471278 16764 471284 16766
rect 471348 16764 471354 16828
rect 416078 16628 416084 16692
rect 416148 16690 416154 16692
rect 511022 16690 511028 16692
rect 416148 16630 511028 16690
rect 416148 16628 416154 16630
rect 511022 16628 511028 16630
rect 511092 16628 511098 16692
rect 357198 7652 357204 7716
rect 357268 7714 357274 7716
rect 534901 7714 534967 7717
rect 357268 7712 534967 7714
rect 357268 7656 534906 7712
rect 534962 7656 534967 7712
rect 357268 7654 534967 7656
rect 357268 7652 357274 7654
rect 534901 7651 534967 7654
rect 359958 7516 359964 7580
rect 360028 7578 360034 7580
rect 541985 7578 542051 7581
rect 360028 7576 542051 7578
rect 360028 7520 541990 7576
rect 542046 7520 542051 7576
rect 360028 7518 542051 7520
rect 360028 7516 360034 7518
rect 541985 7515 542051 7518
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 219157 3906 219223 3909
rect 276013 3906 276079 3909
rect 219157 3904 276079 3906
rect 219157 3848 219162 3904
rect 219218 3848 276018 3904
rect 276074 3848 276079 3904
rect 219157 3846 276079 3848
rect 219157 3843 219223 3846
rect 276013 3843 276079 3846
rect 219801 3770 219867 3773
rect 279509 3770 279575 3773
rect 219801 3768 279575 3770
rect 219801 3712 219806 3768
rect 219862 3712 279514 3768
rect 279570 3712 279575 3768
rect 219801 3710 279575 3712
rect 219801 3707 219867 3710
rect 279509 3707 279575 3710
rect 419942 3708 419948 3772
rect 420012 3770 420018 3772
rect 485221 3770 485287 3773
rect 420012 3768 485287 3770
rect 420012 3712 485226 3768
rect 485282 3712 485287 3768
rect 420012 3710 485287 3712
rect 420012 3708 420018 3710
rect 485221 3707 485287 3710
rect 217133 3634 217199 3637
rect 283097 3634 283163 3637
rect 217133 3632 283163 3634
rect 217133 3576 217138 3632
rect 217194 3576 283102 3632
rect 283158 3576 283163 3632
rect 217133 3574 283163 3576
rect 217133 3571 217199 3574
rect 283097 3571 283163 3574
rect 419758 3572 419764 3636
rect 419828 3634 419834 3636
rect 499389 3634 499455 3637
rect 419828 3632 499455 3634
rect 419828 3576 499394 3632
rect 499450 3576 499455 3632
rect 419828 3574 499455 3576
rect 419828 3572 419834 3574
rect 499389 3571 499455 3574
rect 217225 3498 217291 3501
rect 286593 3498 286659 3501
rect 217225 3496 286659 3498
rect 217225 3440 217230 3496
rect 217286 3440 286598 3496
rect 286654 3440 286659 3496
rect 217225 3438 286659 3440
rect 217225 3435 217291 3438
rect 286593 3435 286659 3438
rect 414749 3498 414815 3501
rect 517145 3498 517211 3501
rect 414749 3496 517211 3498
rect 414749 3440 414754 3496
rect 414810 3440 517150 3496
rect 517206 3440 517211 3496
rect 414749 3438 517211 3440
rect 414749 3435 414815 3438
rect 517145 3435 517211 3438
rect 218881 3362 218947 3365
rect 290181 3362 290247 3365
rect 218881 3360 290247 3362
rect 218881 3304 218886 3360
rect 218942 3304 290186 3360
rect 290242 3304 290247 3360
rect 218881 3302 290247 3304
rect 218881 3299 218947 3302
rect 290181 3299 290247 3302
rect 414933 3362 414999 3365
rect 520733 3362 520799 3365
rect 414933 3360 520799 3362
rect 414933 3304 414938 3360
rect 414994 3304 520738 3360
rect 520794 3304 520799 3360
rect 414933 3302 520799 3304
rect 414933 3299 414999 3302
rect 520733 3299 520799 3302
<< via3 >>
rect 203196 700844 203260 700908
rect 202460 700708 202524 700772
rect 202276 700572 202340 700636
rect 202092 700436 202156 700500
rect 415900 700436 415964 700500
rect 199332 700300 199396 700364
rect 202644 700300 202708 700364
rect 418660 700300 418724 700364
rect 203564 682620 203628 682684
rect 374132 682620 374196 682684
rect 203748 682484 203812 682548
rect 375420 682484 375484 682548
rect 203380 682348 203444 682412
rect 378180 682348 378244 682412
rect 373764 682212 373828 682276
rect 372660 682076 372724 682140
rect 199884 680444 199948 680508
rect 195836 680308 195900 680372
rect 264468 679688 264532 679692
rect 264468 679632 264518 679688
rect 264518 679632 264532 679688
rect 264468 679628 264532 679632
rect 269252 679688 269316 679692
rect 269252 679632 269302 679688
rect 269302 679632 269316 679688
rect 269252 679628 269316 679632
rect 264468 678268 264532 678332
rect 269252 678132 269316 678196
rect 150940 674928 151004 674932
rect 150940 674872 150990 674928
rect 150990 674872 151004 674928
rect 150940 674868 151004 674872
rect 550956 674928 551020 674932
rect 550956 674872 551006 674928
rect 551006 674872 551020 674928
rect 550956 674868 551020 674872
rect 417924 622780 417988 622844
rect 417556 618156 417620 618220
rect 18644 598028 18708 598092
rect 37044 587828 37108 587892
rect 39620 587888 39684 587892
rect 39620 587832 39634 587888
rect 39634 587832 39684 587888
rect 39620 587828 39684 587832
rect 43116 587828 43180 587892
rect 44220 587888 44284 587892
rect 44220 587832 44234 587888
rect 44234 587832 44284 587888
rect 44220 587828 44284 587832
rect 45324 587888 45388 587892
rect 45324 587832 45338 587888
rect 45338 587832 45388 587888
rect 45324 587828 45388 587832
rect 46612 587828 46676 587892
rect 47716 587828 47780 587892
rect 48268 587828 48332 587892
rect 50660 587828 50724 587892
rect 51212 587828 51276 587892
rect 52316 587888 52380 587892
rect 52316 587832 52366 587888
rect 52366 587832 52380 587888
rect 52316 587828 52380 587832
rect 53604 587888 53668 587892
rect 53604 587832 53654 587888
rect 53654 587832 53668 587888
rect 53604 587828 53668 587832
rect 54524 587828 54588 587892
rect 55812 587828 55876 587892
rect 55996 587828 56060 587892
rect 58572 587828 58636 587892
rect 60596 587888 60660 587892
rect 60596 587832 60610 587888
rect 60610 587832 60660 587888
rect 60596 587828 60660 587832
rect 61700 587828 61764 587892
rect 62804 587888 62868 587892
rect 62804 587832 62818 587888
rect 62818 587832 62868 587888
rect 62804 587828 62868 587832
rect 63908 587888 63972 587892
rect 63908 587832 63922 587888
rect 63922 587832 63972 587888
rect 63908 587828 63972 587832
rect 65196 587828 65260 587892
rect 66300 587888 66364 587892
rect 66300 587832 66314 587888
rect 66314 587832 66364 587888
rect 66300 587828 66364 587832
rect 67588 587888 67652 587892
rect 67588 587832 67638 587888
rect 67638 587832 67652 587888
rect 67588 587828 67652 587832
rect 68692 587888 68756 587892
rect 68692 587832 68706 587888
rect 68706 587832 68756 587888
rect 68692 587828 68756 587832
rect 69796 587888 69860 587892
rect 69796 587832 69810 587888
rect 69810 587832 69860 587888
rect 69796 587828 69860 587832
rect 71268 587828 71332 587892
rect 72188 587888 72252 587892
rect 72188 587832 72202 587888
rect 72202 587832 72252 587888
rect 72188 587828 72252 587832
rect 73292 587888 73356 587892
rect 73292 587832 73306 587888
rect 73306 587832 73356 587888
rect 73292 587828 73356 587832
rect 73660 587888 73724 587892
rect 73660 587832 73710 587888
rect 73710 587832 73724 587888
rect 73660 587828 73724 587832
rect 74396 587888 74460 587892
rect 74396 587832 74410 587888
rect 74410 587832 74460 587888
rect 74396 587828 74460 587832
rect 76052 587888 76116 587892
rect 76052 587832 76102 587888
rect 76102 587832 76116 587888
rect 76052 587828 76116 587832
rect 78076 587828 78140 587892
rect 78444 587888 78508 587892
rect 78444 587832 78494 587888
rect 78494 587832 78508 587888
rect 78444 587828 78508 587832
rect 79180 587888 79244 587892
rect 79180 587832 79194 587888
rect 79194 587832 79244 587888
rect 79180 587828 79244 587832
rect 81020 587888 81084 587892
rect 81020 587832 81070 587888
rect 81070 587832 81084 587888
rect 81020 587828 81084 587832
rect 83596 587888 83660 587892
rect 83596 587832 83646 587888
rect 83646 587832 83660 587888
rect 83596 587828 83660 587832
rect 88196 587888 88260 587892
rect 88196 587832 88246 587888
rect 88246 587832 88260 587888
rect 88196 587828 88260 587832
rect 90956 587888 91020 587892
rect 90956 587832 91006 587888
rect 91006 587832 91020 587888
rect 90956 587828 91020 587832
rect 93532 587888 93596 587892
rect 93532 587832 93582 587888
rect 93582 587832 93596 587888
rect 93532 587828 93596 587832
rect 95924 587828 95988 587892
rect 98500 587888 98564 587892
rect 98500 587832 98550 587888
rect 98550 587832 98564 587888
rect 98500 587828 98564 587832
rect 100892 587888 100956 587892
rect 100892 587832 100942 587888
rect 100942 587832 100956 587888
rect 100892 587828 100956 587832
rect 103468 587828 103532 587892
rect 105860 587828 105924 587892
rect 108436 587888 108500 587892
rect 108436 587832 108450 587888
rect 108450 587832 108500 587888
rect 108436 587828 108500 587832
rect 111012 587828 111076 587892
rect 113404 587828 113468 587892
rect 115796 587828 115860 587892
rect 118372 587828 118436 587892
rect 120948 587828 121012 587892
rect 125916 587888 125980 587892
rect 125916 587832 125966 587888
rect 125966 587832 125980 587888
rect 125916 587828 125980 587832
rect 437060 587828 437124 587892
rect 438164 587888 438228 587892
rect 438164 587832 438178 587888
rect 438178 587832 438228 587888
rect 438164 587828 438228 587832
rect 439636 587888 439700 587892
rect 439636 587832 439650 587888
rect 439650 587832 439700 587888
rect 439636 587828 439700 587832
rect 441660 587888 441724 587892
rect 441660 587832 441674 587888
rect 441674 587832 441724 587888
rect 441660 587828 441724 587832
rect 443132 587888 443196 587892
rect 443132 587832 443146 587888
rect 443146 587832 443196 587888
rect 443132 587828 443196 587832
rect 444236 587888 444300 587892
rect 444236 587832 444250 587888
rect 444250 587832 444300 587888
rect 444236 587828 444300 587832
rect 445524 587828 445588 587892
rect 446444 587888 446508 587892
rect 446444 587832 446494 587888
rect 446494 587832 446508 587888
rect 446444 587828 446508 587832
rect 447548 587828 447612 587892
rect 448652 587828 448716 587892
rect 449940 587888 450004 587892
rect 449940 587832 449954 587888
rect 449954 587832 450004 587888
rect 449940 587828 450004 587832
rect 450676 587888 450740 587892
rect 450676 587832 450690 587888
rect 450690 587832 450740 587888
rect 450676 587828 450740 587832
rect 453620 587888 453684 587892
rect 453620 587832 453634 587888
rect 453634 587832 453684 587888
rect 453620 587828 453684 587832
rect 454540 587888 454604 587892
rect 454540 587832 454590 587888
rect 454590 587832 454604 587888
rect 454540 587828 454604 587832
rect 456196 587828 456260 587892
rect 456932 587828 456996 587892
rect 458036 587828 458100 587892
rect 35940 587692 36004 587756
rect 48636 587752 48700 587756
rect 48636 587696 48650 587752
rect 48650 587696 48700 587752
rect 48636 587692 48700 587696
rect 50108 587752 50172 587756
rect 50108 587696 50122 587752
rect 50122 587696 50172 587752
rect 50108 587692 50172 587696
rect 53420 587692 53484 587756
rect 59492 587692 59556 587756
rect 19748 587556 19812 587620
rect 38148 587556 38212 587620
rect 58204 587556 58268 587620
rect 418844 587692 418908 587756
rect 448284 587692 448348 587756
rect 452332 587752 452396 587756
rect 452332 587696 452382 587752
rect 452382 587696 452396 587752
rect 452332 587692 452396 587696
rect 453436 587752 453500 587756
rect 453436 587696 453486 587752
rect 453486 587696 453500 587752
rect 453436 587692 453500 587696
rect 455828 587692 455892 587756
rect 459324 587692 459388 587756
rect 460612 587752 460676 587756
rect 460612 587696 460662 587752
rect 460662 587696 460676 587752
rect 460612 587692 460676 587696
rect 460980 587752 461044 587756
rect 460980 587696 460994 587752
rect 460994 587696 461044 587752
rect 460980 587692 461044 587696
rect 461716 587692 461780 587756
rect 463556 587692 463620 587756
rect 463924 587752 463988 587756
rect 463924 587696 463938 587752
rect 463938 587696 463988 587752
rect 463924 587692 463988 587696
rect 465948 587692 466012 587756
rect 466316 587752 466380 587756
rect 466316 587696 466330 587752
rect 466330 587696 466380 587752
rect 466316 587692 466380 587696
rect 467604 587752 467668 587756
rect 467604 587696 467618 587752
rect 467618 587696 467668 587752
rect 467604 587692 467668 587696
rect 468708 587752 468772 587756
rect 468708 587696 468722 587752
rect 468722 587696 468772 587752
rect 468708 587692 468772 587696
rect 469812 587752 469876 587756
rect 471284 587888 471348 587892
rect 471284 587832 471298 587888
rect 471298 587832 471348 587888
rect 471284 587828 471348 587832
rect 472204 587888 472268 587892
rect 472204 587832 472218 587888
rect 472218 587832 472268 587888
rect 472204 587828 472268 587832
rect 473308 587888 473372 587892
rect 473308 587832 473358 587888
rect 473358 587832 473372 587888
rect 473308 587828 473372 587832
rect 474412 587828 474476 587892
rect 476988 587888 477052 587892
rect 476988 587832 477002 587888
rect 477002 587832 477052 587888
rect 476988 587828 477052 587832
rect 478092 587888 478156 587892
rect 478092 587832 478106 587888
rect 478106 587832 478156 587888
rect 478092 587828 478156 587832
rect 479196 587888 479260 587892
rect 479196 587832 479210 587888
rect 479210 587832 479260 587888
rect 479196 587828 479260 587832
rect 480852 587828 480916 587892
rect 483428 587828 483492 587892
rect 486004 587828 486068 587892
rect 488212 587828 488276 587892
rect 493364 587828 493428 587892
rect 495940 587828 496004 587892
rect 498516 587828 498580 587892
rect 500908 587888 500972 587892
rect 500908 587832 500958 587888
rect 500958 587832 500972 587888
rect 500908 587828 500972 587832
rect 503484 587828 503548 587892
rect 505876 587828 505940 587892
rect 508452 587828 508516 587892
rect 511028 587828 511092 587892
rect 513420 587888 513484 587892
rect 513420 587832 513434 587888
rect 513434 587832 513484 587888
rect 513420 587828 513484 587832
rect 515812 587828 515876 587892
rect 517468 587828 517532 587892
rect 518388 587828 518452 587892
rect 520964 587828 521028 587892
rect 523356 587888 523420 587892
rect 523356 587832 523370 587888
rect 523370 587832 523420 587888
rect 523356 587828 523420 587832
rect 525932 587888 525996 587892
rect 525932 587832 525946 587888
rect 525946 587832 525996 587888
rect 525932 587828 525996 587832
rect 469812 587696 469826 587752
rect 469826 587696 469876 587752
rect 469812 587692 469876 587696
rect 19932 587420 19996 587484
rect 40540 587420 40604 587484
rect 57100 587480 57164 587484
rect 57100 587424 57114 587480
rect 57114 587424 57164 587480
rect 57100 587420 57164 587424
rect 65932 587480 65996 587484
rect 65932 587424 65982 587480
rect 65982 587424 65996 587480
rect 65932 587420 65996 587424
rect 68324 587420 68388 587484
rect 75684 587556 75748 587620
rect 473492 587556 473556 587620
rect 76972 587420 77036 587484
rect 476068 587420 476132 587484
rect 19012 587284 19076 587348
rect 41828 587284 41892 587348
rect 61148 587284 61212 587348
rect 63540 587284 63604 587348
rect 85988 587284 86052 587348
rect 195100 587284 195164 587348
rect 478460 587284 478524 587348
rect 58204 587148 58268 587212
rect 70900 587148 70964 587212
rect 198044 587148 198108 587212
rect 122788 587012 122852 587076
rect 419764 587012 419828 587076
rect 436140 587012 436204 587076
rect 458404 587148 458468 587212
rect 462820 587208 462884 587212
rect 462820 587152 462834 587208
rect 462834 587152 462884 587208
rect 462820 587148 462884 587152
rect 465212 587208 465276 587212
rect 465212 587152 465226 587208
rect 465226 587152 465276 587208
rect 465212 587148 465276 587152
rect 468340 587012 468404 587076
rect 417372 586876 417436 586940
rect 451412 586936 451476 586940
rect 451412 586880 451426 586936
rect 451426 586880 451476 586936
rect 451412 586876 451476 586880
rect 475700 586876 475764 586940
rect 417740 586740 417804 586804
rect 440556 586740 440620 586804
rect 470548 586528 470612 586532
rect 470548 586472 470598 586528
rect 470598 586472 470612 586528
rect 470548 586468 470612 586472
rect 489868 586528 489932 586532
rect 489868 586472 489918 586528
rect 489918 586472 489932 586528
rect 489868 586468 489932 586472
rect 199516 585652 199580 585716
rect 376340 585652 376404 585716
rect 517468 585652 517532 585716
rect 150756 585304 150820 585308
rect 150756 585248 150770 585304
rect 150770 585248 150820 585304
rect 150756 585244 150820 585248
rect 550772 585304 550836 585308
rect 550772 585248 550822 585304
rect 550822 585248 550836 585304
rect 550772 585244 550836 585248
rect 419396 584836 419460 584900
rect 197860 584564 197924 584628
rect 201356 584428 201420 584492
rect 199700 584292 199764 584356
rect 374500 584292 374564 584356
rect 199884 577084 199948 577148
rect 199884 576812 199948 576876
rect 417924 532884 417988 532948
rect 417556 528124 417620 528188
rect 17908 527172 17972 527236
rect 417556 527172 417620 527236
rect 17908 521460 17972 521524
rect 199700 505140 199764 505204
rect 200068 505140 200132 505204
rect 248460 501604 248524 501668
rect 202460 500788 202524 500852
rect 202276 500652 202340 500716
rect 375420 500652 375484 500716
rect 202092 500516 202156 500580
rect 203380 500380 203444 500444
rect 203196 499972 203260 500036
rect 202644 499836 202708 499900
rect 45438 499564 45502 499628
rect 199700 499564 199764 499628
rect 200068 499564 200132 499628
rect 199516 499428 199580 499492
rect 38148 498068 38212 498132
rect 41828 498128 41892 498132
rect 41828 498072 41878 498128
rect 41878 498072 41892 498128
rect 41828 498068 41892 498072
rect 43116 498068 43180 498132
rect 46612 498068 46676 498132
rect 47532 498128 47596 498132
rect 47532 498072 47582 498128
rect 47582 498072 47596 498128
rect 47532 498068 47596 498072
rect 48636 498128 48700 498132
rect 48636 498072 48686 498128
rect 48686 498072 48700 498128
rect 48636 498068 48700 498072
rect 51396 498128 51460 498132
rect 51396 498072 51446 498128
rect 51446 498072 51460 498128
rect 51396 498068 51460 498072
rect 52316 498068 52380 498132
rect 53420 498128 53484 498132
rect 53420 498072 53470 498128
rect 53470 498072 53484 498128
rect 53420 498068 53484 498072
rect 54524 498068 54588 498132
rect 55812 498128 55876 498132
rect 55812 498072 55862 498128
rect 55862 498072 55876 498128
rect 55812 498068 55876 498072
rect 59492 498128 59556 498132
rect 59492 498072 59542 498128
rect 59542 498072 59556 498128
rect 59492 498068 59556 498072
rect 60596 498128 60660 498132
rect 60596 498072 60646 498128
rect 60646 498072 60660 498128
rect 60596 498068 60660 498072
rect 63540 498068 63604 498132
rect 63908 498068 63972 498132
rect 67588 498128 67652 498132
rect 67588 498072 67638 498128
rect 67638 498072 67652 498128
rect 67588 498068 67652 498072
rect 71268 498128 71332 498132
rect 71268 498072 71282 498128
rect 71282 498072 71332 498128
rect 71268 498068 71332 498072
rect 72188 498068 72252 498132
rect 73660 498128 73724 498132
rect 73660 498072 73710 498128
rect 73710 498072 73724 498128
rect 73660 498068 73724 498072
rect 74396 498068 74460 498132
rect 78076 498128 78140 498132
rect 78076 498072 78126 498128
rect 78126 498072 78140 498128
rect 78076 498068 78140 498072
rect 113404 498068 113468 498132
rect 120948 498068 121012 498132
rect 417740 498068 417804 498132
rect 440556 498068 440620 498132
rect 441660 498128 441724 498132
rect 441660 498072 441674 498128
rect 441674 498072 441724 498128
rect 441660 498068 441724 498072
rect 445340 498128 445404 498132
rect 445340 498072 445354 498128
rect 445354 498072 445404 498128
rect 445340 498068 445404 498072
rect 448652 498068 448716 498132
rect 451044 498068 451108 498132
rect 452332 498128 452396 498132
rect 452332 498072 452382 498128
rect 452382 498072 452396 498128
rect 452332 498068 452396 498072
rect 454540 498128 454604 498132
rect 454540 498072 454590 498128
rect 454590 498072 454604 498128
rect 454540 498068 454604 498072
rect 456196 498068 456260 498132
rect 469812 498068 469876 498132
rect 473308 498128 473372 498132
rect 473308 498072 473358 498128
rect 473358 498072 473372 498128
rect 473308 498068 473372 498072
rect 473676 498068 473740 498132
rect 480852 498068 480916 498132
rect 495940 498068 496004 498132
rect 505876 498068 505940 498132
rect 513420 498068 513484 498132
rect 520964 498068 521028 498132
rect 44220 497992 44284 497996
rect 44220 497936 44234 497992
rect 44234 497936 44284 497992
rect 44220 497932 44284 497936
rect 58204 497992 58268 497996
rect 58204 497936 58218 497992
rect 58218 497936 58268 497992
rect 58204 497932 58268 497936
rect 76972 497932 77036 497996
rect 195836 497932 195900 497996
rect 419396 497932 419460 497996
rect 463924 497932 463988 497996
rect 468708 497932 468772 497996
rect 36124 497856 36188 497860
rect 36124 497800 36174 497856
rect 36174 497800 36188 497856
rect 36124 497796 36188 497800
rect 37228 497856 37292 497860
rect 37228 497800 37242 497856
rect 37242 497800 37292 497856
rect 37228 497796 37292 497800
rect 50108 497796 50172 497860
rect 57100 497856 57164 497860
rect 57100 497800 57114 497856
rect 57114 497800 57164 497856
rect 57100 497796 57164 497800
rect 75684 497796 75748 497860
rect 199884 497796 199948 497860
rect 460612 497856 460676 497860
rect 460612 497800 460626 497856
rect 460626 497800 460676 497856
rect 460612 497796 460676 497800
rect 462820 497796 462884 497860
rect 73292 497660 73356 497724
rect 471284 497660 471348 497724
rect 475700 497660 475764 497724
rect 476988 497660 477052 497724
rect 19932 497524 19996 497588
rect 378180 497524 378244 497588
rect 444236 497448 444300 497452
rect 444236 497392 444250 497448
rect 444250 497392 444300 497448
rect 444236 497388 444300 497392
rect 450124 497388 450188 497452
rect 458036 497388 458100 497452
rect 467604 497388 467668 497452
rect 461716 497252 461780 497316
rect 466316 497252 466380 497316
rect 479196 497252 479260 497316
rect 68692 497116 68756 497180
rect 106044 497176 106108 497180
rect 106044 497120 106094 497176
rect 106094 497120 106108 497176
rect 106044 497116 106108 497120
rect 446628 497176 446692 497180
rect 446628 497120 446678 497176
rect 446678 497120 446692 497176
rect 446628 497116 446692 497120
rect 465212 497116 465276 497180
rect 474412 497116 474476 497180
rect 39620 497040 39684 497044
rect 39620 496984 39670 497040
rect 39670 496984 39684 497040
rect 39620 496980 39684 496984
rect 61700 496980 61764 497044
rect 66300 497040 66364 497044
rect 66300 496984 66314 497040
rect 66314 496984 66364 497040
rect 66300 496980 66364 496984
rect 437060 496980 437124 497044
rect 447732 497040 447796 497044
rect 447732 496984 447782 497040
rect 447782 496984 447796 497040
rect 447732 496980 447796 496984
rect 453436 496980 453500 497044
rect 472204 496980 472268 497044
rect 478460 496980 478524 497044
rect 40540 496904 40604 496908
rect 40540 496848 40590 496904
rect 40590 496848 40604 496904
rect 40540 496844 40604 496848
rect 48268 496904 48332 496908
rect 48268 496848 48318 496904
rect 48318 496848 48332 496904
rect 48268 496844 48332 496848
rect 50844 496844 50908 496908
rect 53604 496844 53668 496908
rect 56180 496844 56244 496908
rect 58572 496844 58636 496908
rect 61148 496844 61212 496908
rect 62804 496904 62868 496908
rect 62804 496848 62818 496904
rect 62818 496848 62868 496904
rect 62804 496844 62868 496848
rect 65380 496844 65444 496908
rect 65932 496844 65996 496908
rect 68324 496844 68388 496908
rect 69796 496844 69860 496908
rect 70900 496844 70964 496908
rect 73292 496844 73356 496908
rect 76052 496844 76116 496908
rect 78444 496844 78508 496908
rect 79180 496844 79244 496908
rect 81020 496844 81084 496908
rect 83596 496844 83660 496908
rect 85988 496844 86052 496908
rect 88196 496904 88260 496908
rect 88196 496848 88246 496904
rect 88246 496848 88260 496904
rect 88196 496844 88260 496848
rect 90956 496904 91020 496908
rect 90956 496848 91006 496904
rect 91006 496848 91020 496904
rect 90956 496844 91020 496848
rect 93532 496844 93596 496908
rect 95924 496844 95988 496908
rect 98500 496844 98564 496908
rect 100892 496904 100956 496908
rect 100892 496848 100942 496904
rect 100942 496848 100956 496904
rect 100892 496844 100956 496848
rect 103468 496844 103532 496908
rect 108620 496844 108684 496908
rect 111012 496844 111076 496908
rect 115796 496904 115860 496908
rect 115796 496848 115846 496904
rect 115846 496848 115860 496904
rect 115796 496844 115860 496848
rect 118556 496904 118620 496908
rect 118556 496848 118606 496904
rect 118606 496848 118620 496904
rect 118556 496844 118620 496848
rect 123340 496844 123404 496908
rect 125916 496844 125980 496908
rect 436140 496904 436204 496908
rect 436140 496848 436154 496904
rect 436154 496848 436204 496904
rect 436140 496844 436204 496848
rect 438348 496844 438412 496908
rect 439636 496844 439700 496908
rect 440556 496844 440620 496908
rect 443132 496844 443196 496908
rect 448284 496844 448348 496908
rect 450676 496844 450740 496908
rect 453620 496844 453684 496908
rect 455828 496844 455892 496908
rect 456932 496904 456996 496908
rect 456932 496848 456946 496904
rect 456946 496848 456996 496904
rect 456932 496844 456996 496848
rect 458404 496844 458468 496908
rect 459508 496904 459572 496908
rect 459508 496848 459522 496904
rect 459522 496848 459572 496904
rect 459508 496844 459572 496848
rect 460980 496904 461044 496908
rect 460980 496848 460994 496904
rect 460994 496848 461044 496904
rect 460980 496844 461044 496848
rect 463556 496844 463620 496908
rect 465948 496844 466012 496908
rect 468340 496844 468404 496908
rect 470916 496844 470980 496908
rect 476068 496904 476132 496908
rect 476068 496848 476118 496904
rect 476118 496848 476132 496904
rect 476068 496844 476132 496848
rect 478092 496844 478156 496908
rect 483428 496844 483492 496908
rect 486004 496844 486068 496908
rect 488212 496844 488276 496908
rect 490972 496844 491036 496908
rect 493364 496844 493428 496908
rect 498516 496844 498580 496908
rect 500908 496904 500972 496908
rect 500908 496848 500958 496904
rect 500958 496848 500972 496904
rect 500908 496844 500972 496848
rect 503484 496844 503548 496908
rect 508452 496844 508516 496908
rect 511028 496844 511092 496908
rect 515812 496844 515876 496908
rect 518388 496844 518452 496908
rect 523356 496844 523420 496908
rect 525932 496844 525996 496908
rect 419764 496708 419828 496772
rect 18644 496028 18708 496092
rect 374132 494940 374196 495004
rect 372660 494804 372724 494868
rect 19012 494668 19076 494732
rect 373764 494668 373828 494732
rect 417372 493988 417436 494052
rect 418844 493308 418908 493372
rect 19748 491132 19812 491196
rect 418660 480796 418724 480860
rect 195100 475356 195164 475420
rect 199332 468420 199396 468484
rect 203564 466108 203628 466172
rect 198044 465836 198108 465900
rect 192708 463660 192772 463724
rect 417372 463720 417436 463724
rect 417372 463664 417422 463720
rect 417422 463664 417436 463720
rect 417372 463660 417436 463664
rect 199884 461620 199948 461684
rect 201356 461484 201420 461548
rect 192156 461348 192220 461412
rect 197860 460124 197924 460188
rect 188476 458900 188540 458964
rect 415900 457404 415964 457468
rect 186820 457268 186884 457332
rect 184060 457132 184124 457196
rect 19196 456860 19260 456924
rect 187004 456044 187068 456108
rect 187188 455908 187252 455972
rect 184244 455772 184308 455836
rect 190316 454684 190380 454748
rect 188292 454548 188356 454612
rect 191052 454412 191116 454476
rect 18460 454276 18524 454340
rect 414612 454276 414676 454340
rect 185164 453188 185228 453252
rect 192524 453052 192588 453116
rect 418108 453052 418172 453116
rect 248460 452508 248524 452572
rect 374500 452508 374564 452572
rect 376340 452508 376404 452572
rect 418660 452372 418724 452436
rect 418844 452236 418908 452300
rect 203748 452100 203812 452164
rect 415900 451828 415964 451892
rect 419028 451692 419092 451756
rect 188844 451480 188908 451484
rect 188844 451424 188894 451480
rect 188894 451424 188908 451480
rect 188844 451420 188908 451424
rect 188660 451284 188724 451348
rect 191604 451284 191668 451348
rect 417740 450876 417804 450940
rect 191236 450740 191300 450804
rect 192340 450604 192404 450668
rect 191420 450468 191484 450532
rect 187372 450332 187436 450396
rect 193812 450196 193876 450260
rect 416084 449788 416148 449852
rect 190132 449652 190196 449716
rect 389220 449652 389284 449716
rect 193996 449304 194060 449308
rect 193996 449248 194046 449304
rect 194046 449248 194060 449304
rect 193996 449244 194060 449248
rect 417556 449108 417620 449172
rect 192340 395932 192404 395996
rect 192340 394708 192404 394772
rect 192156 369820 192220 369884
rect 191788 369200 191852 369204
rect 191788 369144 191838 369200
rect 191838 369144 191852 369200
rect 191788 369140 191852 369144
rect 190132 249052 190196 249116
rect 357204 247148 357268 247212
rect 359964 247012 360028 247076
rect 150940 196072 151004 196076
rect 150940 196016 150990 196072
rect 150990 196016 151004 196072
rect 150940 196012 151004 196016
rect 550956 196072 551020 196076
rect 550956 196016 551006 196072
rect 551006 196016 551020 196072
rect 550956 196012 551020 196016
rect 193996 193972 194060 194036
rect 193812 193836 193876 193900
rect 417188 145964 417252 146028
rect 417740 145964 417804 146028
rect 417740 142700 417804 142764
rect 417556 138212 417620 138276
rect 417924 138212 417988 138276
rect 419764 111148 419828 111212
rect 419948 111012 420012 111076
rect 451286 109848 451350 109852
rect 451286 109792 451334 109848
rect 451334 109792 451350 109848
rect 451286 109788 451350 109792
rect 480934 109848 480998 109852
rect 480934 109792 480958 109848
rect 480958 109792 480998 109848
rect 480934 109788 480998 109792
rect 483518 109848 483582 109852
rect 483518 109792 483534 109848
rect 483534 109792 483582 109848
rect 483518 109788 483582 109792
rect 485966 109848 486030 109852
rect 485966 109792 486018 109848
rect 486018 109792 486030 109848
rect 485966 109788 486030 109792
rect 488278 109848 488342 109852
rect 488278 109792 488318 109848
rect 488318 109792 488342 109848
rect 488278 109788 488342 109792
rect 490998 109848 491062 109852
rect 490998 109792 491022 109848
rect 491022 109792 491062 109848
rect 490998 109788 491062 109792
rect 476068 109712 476132 109716
rect 476068 109656 476118 109712
rect 476118 109656 476132 109712
rect 476068 109652 476132 109656
rect 493446 109712 493510 109716
rect 493446 109656 493470 109712
rect 493470 109656 493510 109712
rect 493446 109652 493510 109656
rect 495894 109712 495958 109716
rect 495894 109656 495898 109712
rect 495898 109656 495954 109712
rect 495954 109656 495958 109712
rect 495894 109652 495958 109656
rect 498478 109712 498542 109716
rect 498478 109656 498530 109712
rect 498530 109656 498542 109712
rect 498478 109652 498542 109656
rect 50742 109576 50806 109580
rect 50742 109520 50802 109576
rect 50802 109520 50806 109576
rect 50742 109516 50806 109520
rect 56046 109576 56110 109580
rect 56046 109520 56102 109576
rect 56102 109520 56110 109576
rect 56046 109516 56110 109520
rect 61078 109576 61142 109580
rect 61078 109520 61106 109576
rect 61106 109520 61142 109576
rect 61078 109516 61142 109520
rect 105958 109576 106022 109580
rect 105958 109520 106002 109576
rect 106002 109520 106022 109576
rect 105958 109516 106022 109520
rect 108542 109576 108606 109580
rect 108542 109520 108578 109576
rect 108578 109520 108606 109576
rect 108542 109516 108606 109520
rect 456998 109576 457062 109580
rect 456998 109520 457038 109576
rect 457038 109520 457062 109576
rect 456998 109516 457062 109520
rect 461078 109516 461142 109580
rect 505958 109576 506022 109580
rect 505958 109520 505982 109576
rect 505982 109520 506022 109576
rect 505958 109516 506022 109520
rect 508542 109576 508606 109580
rect 508542 109520 508558 109576
rect 508558 109520 508606 109576
rect 508542 109516 508606 109520
rect 515886 109576 515950 109580
rect 515886 109520 515918 109576
rect 515918 109520 515950 109576
rect 515886 109516 515950 109520
rect 518470 109576 518534 109580
rect 518470 109520 518494 109576
rect 518494 109520 518534 109576
rect 518470 109516 518534 109520
rect 468340 109108 468404 109172
rect 48268 109032 48332 109036
rect 48268 108976 48318 109032
rect 48318 108976 48332 109032
rect 48268 108972 48332 108976
rect 68324 109032 68388 109036
rect 68324 108976 68374 109032
rect 68374 108976 68388 109032
rect 68324 108972 68388 108976
rect 100892 109032 100956 109036
rect 100892 108976 100942 109032
rect 100942 108976 100956 109032
rect 100892 108972 100956 108976
rect 111012 109032 111076 109036
rect 111012 108976 111062 109032
rect 111062 108976 111076 109032
rect 111012 108972 111076 108976
rect 113404 109032 113468 109036
rect 113404 108976 113454 109032
rect 113454 108976 113468 109032
rect 113404 108972 113468 108976
rect 125916 108972 125980 109036
rect 389220 108972 389284 109036
rect 470916 108972 470980 109036
rect 500908 109032 500972 109036
rect 500908 108976 500958 109032
rect 500958 108976 500972 109032
rect 500908 108972 500972 108976
rect 503484 109032 503548 109036
rect 503484 108976 503498 109032
rect 503498 108976 503548 109032
rect 503484 108972 503548 108976
rect 513420 109032 513484 109036
rect 513420 108976 513434 109032
rect 513434 108976 513484 109032
rect 513420 108972 513484 108976
rect 520964 109032 521028 109036
rect 520964 108976 520978 109032
rect 520978 108976 521028 109032
rect 520964 108972 521028 108976
rect 523356 109032 523420 109036
rect 523356 108976 523370 109032
rect 523370 108976 523420 109032
rect 523356 108972 523420 108976
rect 525932 109032 525996 109036
rect 525932 108976 525946 109032
rect 525946 108976 525996 109032
rect 525932 108972 525996 108976
rect 65932 108836 65996 108900
rect 188476 108836 188540 108900
rect 465948 108836 466012 108900
rect 53604 108760 53668 108764
rect 53604 108704 53654 108760
rect 53654 108704 53668 108760
rect 53604 108700 53668 108704
rect 90956 108700 91020 108764
rect 186820 108700 186884 108764
rect 95924 108564 95988 108628
rect 187188 108564 187252 108628
rect 118556 108428 118620 108492
rect 184244 108428 184308 108492
rect 458036 108488 458100 108492
rect 458036 108432 458050 108488
rect 458050 108432 458100 108488
rect 458036 108428 458100 108432
rect 19932 107476 19996 107540
rect 35940 107536 36004 107540
rect 35940 107480 35954 107536
rect 35954 107480 36004 107536
rect 35940 107476 36004 107480
rect 37044 107476 37108 107540
rect 38148 107536 38212 107540
rect 38148 107480 38162 107536
rect 38162 107480 38212 107536
rect 38148 107476 38212 107480
rect 39620 107536 39684 107540
rect 39620 107480 39634 107536
rect 39634 107480 39684 107536
rect 39620 107476 39684 107480
rect 40540 107536 40604 107540
rect 40540 107480 40554 107536
rect 40554 107480 40604 107536
rect 40540 107476 40604 107480
rect 43116 107536 43180 107540
rect 43116 107480 43166 107536
rect 43166 107480 43180 107536
rect 43116 107476 43180 107480
rect 44220 107536 44284 107540
rect 44220 107480 44270 107536
rect 44270 107480 44284 107536
rect 44220 107476 44284 107480
rect 45324 107536 45388 107540
rect 45324 107480 45374 107536
rect 45374 107480 45388 107536
rect 45324 107476 45388 107480
rect 46612 107536 46676 107540
rect 46612 107480 46626 107536
rect 46626 107480 46676 107536
rect 46612 107476 46676 107480
rect 47532 107536 47596 107540
rect 47532 107480 47582 107536
rect 47582 107480 47596 107536
rect 47532 107476 47596 107480
rect 48636 107476 48700 107540
rect 50108 107536 50172 107540
rect 50108 107480 50158 107536
rect 50158 107480 50172 107536
rect 50108 107476 50172 107480
rect 51212 107536 51276 107540
rect 51212 107480 51262 107536
rect 51262 107480 51276 107536
rect 51212 107476 51276 107480
rect 52316 107536 52380 107540
rect 52316 107480 52366 107536
rect 52366 107480 52380 107536
rect 52316 107476 52380 107480
rect 53420 107536 53484 107540
rect 53420 107480 53470 107536
rect 53470 107480 53484 107536
rect 53420 107476 53484 107480
rect 59492 107476 59556 107540
rect 60596 107536 60660 107540
rect 60596 107480 60610 107536
rect 60610 107480 60660 107536
rect 60596 107476 60660 107480
rect 61700 107536 61764 107540
rect 61700 107480 61714 107536
rect 61714 107480 61764 107536
rect 61700 107476 61764 107480
rect 62804 107476 62868 107540
rect 63540 107536 63604 107540
rect 63540 107480 63590 107536
rect 63590 107480 63604 107536
rect 63540 107476 63604 107480
rect 63908 107536 63972 107540
rect 63908 107480 63922 107536
rect 63922 107480 63972 107536
rect 63908 107476 63972 107480
rect 65196 107536 65260 107540
rect 65196 107480 65210 107536
rect 65210 107480 65260 107536
rect 65196 107476 65260 107480
rect 66300 107536 66364 107540
rect 66300 107480 66314 107536
rect 66314 107480 66364 107536
rect 66300 107476 66364 107480
rect 67588 107536 67652 107540
rect 67588 107480 67638 107536
rect 67638 107480 67652 107536
rect 67588 107476 67652 107480
rect 68692 107536 68756 107540
rect 68692 107480 68706 107536
rect 68706 107480 68756 107536
rect 68692 107476 68756 107480
rect 69796 107536 69860 107540
rect 69796 107480 69810 107536
rect 69810 107480 69860 107536
rect 69796 107476 69860 107480
rect 71268 107536 71332 107540
rect 71268 107480 71282 107536
rect 71282 107480 71332 107536
rect 71268 107476 71332 107480
rect 72188 107536 72252 107540
rect 72188 107480 72202 107536
rect 72202 107480 72252 107536
rect 72188 107476 72252 107480
rect 73292 107536 73356 107540
rect 73292 107480 73306 107536
rect 73306 107480 73356 107536
rect 73292 107476 73356 107480
rect 73660 107536 73724 107540
rect 73660 107480 73710 107536
rect 73710 107480 73724 107536
rect 73660 107476 73724 107480
rect 74396 107536 74460 107540
rect 74396 107480 74410 107536
rect 74410 107480 74460 107536
rect 74396 107476 74460 107480
rect 75684 107536 75748 107540
rect 75684 107480 75698 107536
rect 75698 107480 75748 107536
rect 75684 107476 75748 107480
rect 76052 107536 76116 107540
rect 76052 107480 76102 107536
rect 76102 107480 76116 107536
rect 76052 107476 76116 107480
rect 78076 107476 78140 107540
rect 78444 107536 78508 107540
rect 78444 107480 78494 107536
rect 78494 107480 78508 107536
rect 78444 107476 78508 107480
rect 79180 107536 79244 107540
rect 79180 107480 79194 107536
rect 79194 107480 79244 107536
rect 79180 107476 79244 107480
rect 85988 107536 86052 107540
rect 85988 107480 86038 107536
rect 86038 107480 86052 107536
rect 85988 107476 86052 107480
rect 88196 107536 88260 107540
rect 88196 107480 88246 107536
rect 88246 107480 88260 107536
rect 88196 107476 88260 107480
rect 93532 107536 93596 107540
rect 93532 107480 93582 107536
rect 93582 107480 93596 107536
rect 93532 107476 93596 107480
rect 98500 107536 98564 107540
rect 98500 107480 98550 107536
rect 98550 107480 98564 107536
rect 98500 107476 98564 107480
rect 120948 107536 121012 107540
rect 120948 107480 120998 107536
rect 120998 107480 121012 107536
rect 120948 107476 121012 107480
rect 123340 107536 123404 107540
rect 123340 107480 123390 107536
rect 123390 107480 123404 107536
rect 123340 107476 123404 107480
rect 417372 107476 417436 107540
rect 436140 107536 436204 107540
rect 436140 107480 436154 107536
rect 436154 107480 436204 107536
rect 436140 107476 436204 107480
rect 437060 107536 437124 107540
rect 437060 107480 437074 107536
rect 437074 107480 437124 107536
rect 437060 107476 437124 107480
rect 438164 107536 438228 107540
rect 438164 107480 438178 107536
rect 438178 107480 438228 107536
rect 438164 107476 438228 107480
rect 439636 107536 439700 107540
rect 439636 107480 439650 107536
rect 439650 107480 439700 107536
rect 439636 107476 439700 107480
rect 440556 107536 440620 107540
rect 440556 107480 440570 107536
rect 440570 107480 440620 107536
rect 440556 107476 440620 107480
rect 441660 107536 441724 107540
rect 441660 107480 441674 107536
rect 441674 107480 441724 107536
rect 441660 107476 441724 107480
rect 443132 107536 443196 107540
rect 443132 107480 443146 107536
rect 443146 107480 443196 107536
rect 443132 107476 443196 107480
rect 444236 107536 444300 107540
rect 444236 107480 444250 107536
rect 444250 107480 444300 107536
rect 444236 107476 444300 107480
rect 445524 107476 445588 107540
rect 446444 107536 446508 107540
rect 446444 107480 446458 107536
rect 446458 107480 446508 107536
rect 446444 107476 446508 107480
rect 447548 107476 447612 107540
rect 448652 107476 448716 107540
rect 450124 107476 450188 107540
rect 450676 107536 450740 107540
rect 450676 107480 450690 107536
rect 450690 107480 450740 107536
rect 450676 107476 450740 107480
rect 452332 107476 452396 107540
rect 453620 107536 453684 107540
rect 453620 107480 453634 107536
rect 453634 107480 453684 107536
rect 453620 107476 453684 107480
rect 454540 107536 454604 107540
rect 454540 107480 454590 107536
rect 454590 107480 454604 107536
rect 454540 107476 454604 107480
rect 455828 107536 455892 107540
rect 455828 107480 455842 107536
rect 455842 107480 455892 107536
rect 455828 107476 455892 107480
rect 456012 107536 456076 107540
rect 456012 107480 456026 107536
rect 456026 107480 456076 107536
rect 456012 107476 456076 107480
rect 458404 107536 458468 107540
rect 458404 107480 458418 107536
rect 458418 107480 458468 107536
rect 458404 107476 458468 107480
rect 459508 107536 459572 107540
rect 459508 107480 459522 107536
rect 459522 107480 459572 107536
rect 459508 107476 459572 107480
rect 460612 107536 460676 107540
rect 460612 107480 460662 107536
rect 460662 107480 460676 107536
rect 460612 107476 460676 107480
rect 461716 107536 461780 107540
rect 461716 107480 461730 107536
rect 461730 107480 461780 107536
rect 461716 107476 461780 107480
rect 462820 107536 462884 107540
rect 462820 107480 462834 107536
rect 462834 107480 462884 107536
rect 462820 107476 462884 107480
rect 463924 107536 463988 107540
rect 463924 107480 463938 107536
rect 463938 107480 463988 107536
rect 463924 107476 463988 107480
rect 465212 107536 465276 107540
rect 465212 107480 465226 107536
rect 465226 107480 465276 107536
rect 465212 107476 465276 107480
rect 466316 107476 466380 107540
rect 467604 107476 467668 107540
rect 468708 107536 468772 107540
rect 468708 107480 468722 107536
rect 468722 107480 468772 107536
rect 468708 107476 468772 107480
rect 469812 107536 469876 107540
rect 469812 107480 469826 107536
rect 469826 107480 469876 107536
rect 469812 107476 469876 107480
rect 471284 107476 471348 107540
rect 472204 107476 472268 107540
rect 473308 107536 473372 107540
rect 473308 107480 473358 107536
rect 473358 107480 473372 107536
rect 473308 107476 473372 107480
rect 474412 107536 474476 107540
rect 474412 107480 474426 107536
rect 474426 107480 474476 107536
rect 474412 107476 474476 107480
rect 475700 107536 475764 107540
rect 475700 107480 475714 107536
rect 475714 107480 475764 107536
rect 475700 107476 475764 107480
rect 478092 107536 478156 107540
rect 478092 107480 478106 107536
rect 478106 107480 478156 107536
rect 478092 107476 478156 107480
rect 479196 107536 479260 107540
rect 479196 107480 479210 107536
rect 479210 107480 479260 107536
rect 479196 107476 479260 107480
rect 19012 107340 19076 107404
rect 41828 107340 41892 107404
rect 57100 107340 57164 107404
rect 70900 107340 70964 107404
rect 191236 107340 191300 107404
rect 463556 107340 463620 107404
rect 58020 107204 58084 107268
rect 76972 107204 77036 107268
rect 81020 107204 81084 107268
rect 187372 107204 187436 107268
rect 478460 107204 478524 107268
rect 54524 107068 54588 107132
rect 55812 107128 55876 107132
rect 55812 107072 55826 107128
rect 55826 107072 55876 107128
rect 55812 107068 55876 107072
rect 83596 107068 83660 107132
rect 187004 107068 187068 107132
rect 448284 107068 448348 107132
rect 453436 107068 453500 107132
rect 476988 107068 477052 107132
rect 103468 106932 103532 106996
rect 191420 106932 191484 106996
rect 419028 106932 419092 106996
rect 473492 106932 473556 106996
rect 115796 106796 115860 106860
rect 184060 106796 184124 106860
rect 58572 106660 58636 106724
rect 511028 106660 511092 106724
rect 57100 106312 57164 106316
rect 57100 106256 57114 106312
rect 57114 106256 57164 106312
rect 57100 106252 57164 106256
rect 350948 106116 351012 106180
rect 191604 105708 191668 105772
rect 188844 105572 188908 105636
rect 188660 105436 188724 105500
rect 150756 105360 150820 105364
rect 150756 105304 150806 105360
rect 150806 105304 150820 105360
rect 150756 105300 150820 105304
rect 550772 105360 550836 105364
rect 550772 105304 550786 105360
rect 550786 105304 550836 105360
rect 550772 105300 550836 105304
rect 18460 96596 18524 96660
rect 417188 55932 417252 55996
rect 417740 52804 417804 52868
rect 417924 48180 417988 48244
rect 190316 29956 190380 30020
rect 19196 28052 19260 28116
rect 460670 19816 460734 19820
rect 460670 19760 460718 19816
rect 460718 19760 460734 19816
rect 460670 19756 460734 19760
rect 488278 19816 488342 19820
rect 488278 19760 488318 19816
rect 488318 19760 488342 19816
rect 488278 19756 488342 19760
rect 447614 19680 447678 19684
rect 447614 19624 447654 19680
rect 447654 19624 447678 19680
rect 447614 19620 447678 19624
rect 448702 19680 448766 19684
rect 448702 19624 448758 19680
rect 448758 19624 448766 19680
rect 448702 19620 448766 19624
rect 450062 19680 450126 19684
rect 450062 19624 450082 19680
rect 450082 19624 450126 19680
rect 450062 19620 450126 19624
rect 455910 19680 455974 19684
rect 455910 19624 455970 19680
rect 455970 19624 455974 19680
rect 455910 19620 455974 19624
rect 473318 19680 473382 19684
rect 473318 19624 473358 19680
rect 473358 19624 473382 19680
rect 473318 19620 473382 19624
rect 490998 19680 491062 19684
rect 490998 19624 491022 19680
rect 491022 19624 491062 19680
rect 490998 19620 491062 19624
rect 493446 19680 493510 19684
rect 493446 19624 493470 19680
rect 493470 19624 493510 19680
rect 493446 19620 493510 19624
rect 52374 19544 52438 19548
rect 52374 19488 52422 19544
rect 52422 19488 52438 19544
rect 52374 19484 52438 19488
rect 53462 19544 53526 19548
rect 53462 19488 53470 19544
rect 53470 19488 53526 19544
rect 53462 19484 53526 19488
rect 55910 19544 55974 19548
rect 55910 19488 55954 19544
rect 55954 19488 55974 19544
rect 55910 19484 55974 19488
rect 285966 19544 286030 19548
rect 285966 19488 286010 19544
rect 286010 19488 286030 19544
rect 285966 19484 286030 19488
rect 461078 19484 461142 19548
rect 468286 19544 468350 19548
rect 468286 19488 468298 19544
rect 468298 19488 468350 19544
rect 468286 19484 468350 19488
rect 485966 19484 486030 19548
rect 495894 19544 495958 19548
rect 495894 19488 495898 19544
rect 495898 19488 495954 19544
rect 495954 19488 495958 19544
rect 495894 19484 495958 19488
rect 500926 19544 500990 19548
rect 500926 19488 500958 19544
rect 500958 19488 500990 19544
rect 500926 19484 500990 19488
rect 503510 19544 503574 19548
rect 503510 19488 503534 19544
rect 503534 19488 503574 19544
rect 503510 19484 503574 19488
rect 95924 19272 95988 19276
rect 95924 19216 95974 19272
rect 95974 19216 95988 19272
rect 95924 19212 95988 19216
rect 100892 19272 100956 19276
rect 100892 19216 100942 19272
rect 100942 19216 100956 19272
rect 100892 19212 100956 19216
rect 103652 19272 103716 19276
rect 103652 19216 103702 19272
rect 103702 19216 103716 19272
rect 103652 19212 103716 19216
rect 118556 19212 118620 19276
rect 185164 19212 185228 19276
rect 240548 19212 240612 19276
rect 244228 19272 244292 19276
rect 244228 19216 244278 19272
rect 244278 19216 244292 19272
rect 244228 19212 244292 19216
rect 245332 19272 245396 19276
rect 245332 19216 245346 19272
rect 245346 19216 245396 19272
rect 245332 19212 245396 19216
rect 246436 19272 246500 19276
rect 246436 19216 246450 19272
rect 246450 19216 246500 19272
rect 246436 19212 246500 19216
rect 415900 19212 415964 19276
rect 498516 19272 498580 19276
rect 498516 19216 498530 19272
rect 498530 19216 498580 19272
rect 498516 19212 498580 19216
rect 520964 19212 521028 19276
rect 85988 19136 86052 19140
rect 85988 19080 86038 19136
rect 86038 19080 86052 19136
rect 85988 19076 86052 19080
rect 90956 19136 91020 19140
rect 90956 19080 91006 19136
rect 91006 19080 91020 19136
rect 90956 19076 91020 19080
rect 120948 19076 121012 19140
rect 239628 19076 239692 19140
rect 248276 19136 248340 19140
rect 248276 19080 248290 19136
rect 248290 19080 248340 19136
rect 248276 19076 248340 19080
rect 250116 19136 250180 19140
rect 250116 19080 250130 19136
rect 250130 19080 250180 19136
rect 250116 19076 250180 19080
rect 418108 19076 418172 19140
rect 418844 19076 418908 19140
rect 518388 19076 518452 19140
rect 76052 19000 76116 19004
rect 76052 18944 76102 19000
rect 76102 18944 76116 19000
rect 76052 18940 76116 18944
rect 81020 19000 81084 19004
rect 81020 18944 81070 19000
rect 81070 18944 81084 19000
rect 81020 18940 81084 18944
rect 241652 18940 241716 19004
rect 247540 19000 247604 19004
rect 247540 18944 247554 19000
rect 247554 18944 247604 19000
rect 247540 18940 247604 18944
rect 250668 19000 250732 19004
rect 250668 18944 250682 19000
rect 250682 18944 250732 19000
rect 250668 18940 250732 18944
rect 418660 18940 418724 19004
rect 513420 18940 513484 19004
rect 515812 19000 515876 19004
rect 515812 18944 515826 19000
rect 515826 18944 515876 19000
rect 515812 18940 515876 18944
rect 55996 18864 56060 18868
rect 55996 18808 56046 18864
rect 56046 18808 56060 18864
rect 55996 18804 56060 18808
rect 58204 18864 58268 18868
rect 58204 18808 58218 18864
rect 58218 18808 58268 18864
rect 58204 18804 58268 18808
rect 73660 18864 73724 18868
rect 73660 18808 73710 18864
rect 73710 18808 73724 18864
rect 73660 18804 73724 18808
rect 238156 18804 238220 18868
rect 252324 18864 252388 18868
rect 252324 18808 252338 18864
rect 252338 18808 252388 18864
rect 252324 18804 252388 18808
rect 253612 18864 253676 18868
rect 253612 18808 253626 18864
rect 253626 18808 253676 18864
rect 253612 18804 253676 18808
rect 465948 18804 466012 18868
rect 470916 18864 470980 18868
rect 470916 18808 470930 18864
rect 470930 18808 470980 18864
rect 470916 18804 470980 18808
rect 505876 18864 505940 18868
rect 505876 18808 505890 18864
rect 505890 18808 505940 18864
rect 505876 18804 505940 18808
rect 508452 18864 508516 18868
rect 508452 18808 508466 18864
rect 508466 18808 508516 18864
rect 508452 18804 508516 18808
rect 50844 18728 50908 18732
rect 50844 18672 50894 18728
rect 50894 18672 50908 18728
rect 50844 18668 50908 18672
rect 53604 18728 53668 18732
rect 53604 18672 53654 18728
rect 53654 18672 53668 18728
rect 53604 18668 53668 18672
rect 237052 18668 237116 18732
rect 256004 18728 256068 18732
rect 256004 18672 256018 18728
rect 256018 18672 256068 18728
rect 256004 18668 256068 18672
rect 258396 18728 258460 18732
rect 258396 18672 258410 18728
rect 258410 18672 258460 18728
rect 258396 18668 258460 18672
rect 523356 18728 523420 18732
rect 523356 18672 523370 18728
rect 523370 18672 523420 18728
rect 106044 18592 106108 18596
rect 106044 18536 106094 18592
rect 106094 18536 106108 18592
rect 106044 18532 106108 18536
rect 108620 18592 108684 18596
rect 108620 18536 108670 18592
rect 108670 18536 108684 18592
rect 108620 18532 108684 18536
rect 235948 18592 236012 18596
rect 235948 18536 235998 18592
rect 235998 18536 236012 18592
rect 235948 18532 236012 18536
rect 243124 18592 243188 18596
rect 243124 18536 243138 18592
rect 243138 18536 243188 18592
rect 243124 18532 243188 18536
rect 523356 18668 523420 18672
rect 525932 18728 525996 18732
rect 525932 18672 525946 18728
rect 525946 18672 525996 18728
rect 525932 18668 525996 18672
rect 463556 18532 463620 18596
rect 113404 18456 113468 18460
rect 113404 18400 113454 18456
rect 113454 18400 113468 18456
rect 113404 18396 113468 18400
rect 41644 18124 41708 18188
rect 45324 18124 45388 18188
rect 74396 18124 74460 18188
rect 37044 17852 37108 17916
rect 19012 17716 19076 17780
rect 43116 17912 43180 17916
rect 43116 17856 43130 17912
rect 43130 17856 43180 17912
rect 43116 17852 43180 17856
rect 44220 17912 44284 17916
rect 44220 17856 44234 17912
rect 44234 17856 44284 17912
rect 44220 17852 44284 17856
rect 46612 17912 46676 17916
rect 46612 17856 46662 17912
rect 46662 17856 46676 17912
rect 46612 17852 46676 17856
rect 47532 17912 47596 17916
rect 47532 17856 47582 17912
rect 47582 17856 47596 17912
rect 47532 17852 47596 17856
rect 48636 17912 48700 17916
rect 48636 17856 48686 17912
rect 48686 17856 48700 17912
rect 48636 17852 48700 17856
rect 50108 17912 50172 17916
rect 50108 17856 50158 17912
rect 50158 17856 50172 17912
rect 50108 17852 50172 17856
rect 51396 17912 51460 17916
rect 51396 17856 51446 17912
rect 51446 17856 51460 17912
rect 51396 17852 51460 17856
rect 59492 17912 59556 17916
rect 59492 17856 59542 17912
rect 59542 17856 59556 17912
rect 59492 17852 59556 17856
rect 60596 17852 60660 17916
rect 61148 17852 61212 17916
rect 63540 17852 63604 17916
rect 65932 17852 65996 17916
rect 68692 17852 68756 17916
rect 72188 17852 72252 17916
rect 458404 18048 458468 18052
rect 458404 17992 458418 18048
rect 458418 17992 458468 18048
rect 458404 17988 458468 17992
rect 78444 17852 78508 17916
rect 125916 17912 125980 17916
rect 125916 17856 125966 17912
rect 125966 17856 125980 17912
rect 125916 17852 125980 17856
rect 48268 17716 48332 17780
rect 192340 17716 192404 17780
rect 268332 17852 268396 17916
rect 273484 17852 273548 17916
rect 277164 17852 277228 17916
rect 280844 17852 280908 17916
rect 436140 17912 436204 17916
rect 436140 17856 436154 17912
rect 436154 17856 436204 17912
rect 436140 17852 436204 17856
rect 437060 17852 437124 17916
rect 438348 17852 438412 17916
rect 439636 17852 439700 17916
rect 440556 17852 440620 17916
rect 442028 17852 442092 17916
rect 443132 17912 443196 17916
rect 443132 17856 443146 17912
rect 443146 17856 443196 17912
rect 443132 17852 443196 17856
rect 444236 17912 444300 17916
rect 444236 17856 444286 17912
rect 444286 17856 444300 17912
rect 444236 17852 444300 17856
rect 445708 17912 445772 17916
rect 445708 17856 445722 17912
rect 445722 17856 445772 17912
rect 445708 17852 445772 17856
rect 446444 17912 446508 17916
rect 446444 17856 446494 17912
rect 446494 17856 446508 17912
rect 446444 17852 446508 17856
rect 448284 17852 448348 17916
rect 450676 17852 450740 17916
rect 451412 17852 451476 17916
rect 452332 17912 452396 17916
rect 452332 17856 452346 17912
rect 452346 17856 452396 17912
rect 452332 17852 452396 17856
rect 453436 17912 453500 17916
rect 453436 17856 453486 17912
rect 453486 17856 453500 17912
rect 453436 17852 453500 17856
rect 454540 17852 454604 17916
rect 456012 17852 456076 17916
rect 457116 17852 457180 17916
rect 458036 17912 458100 17916
rect 458036 17856 458086 17912
rect 458086 17856 458100 17912
rect 458036 17852 458100 17856
rect 459324 17852 459388 17916
rect 461716 17852 461780 17916
rect 462820 17852 462884 17916
rect 463924 17852 463988 17916
rect 466316 17852 466380 17916
rect 467604 17852 467668 17916
rect 468708 17852 468772 17916
rect 474412 17852 474476 17916
rect 476988 17852 477052 17916
rect 479196 17852 479260 17916
rect 263548 17776 263612 17780
rect 263548 17720 263598 17776
rect 263598 17720 263612 17776
rect 263548 17716 263612 17720
rect 265940 17716 266004 17780
rect 473308 17716 473372 17780
rect 480668 17716 480732 17780
rect 40540 17580 40604 17644
rect 54524 17580 54588 17644
rect 68324 17580 68388 17644
rect 71268 17580 71332 17644
rect 83596 17580 83660 17644
rect 115796 17580 115860 17644
rect 188292 17580 188356 17644
rect 192524 17580 192588 17644
rect 254532 17580 254596 17644
rect 260604 17580 260668 17644
rect 260972 17580 261036 17644
rect 270908 17580 270972 17644
rect 483428 17580 483492 17644
rect 38516 17444 38580 17508
rect 58204 17444 58268 17508
rect 76972 17444 77036 17508
rect 79180 17444 79244 17508
rect 88196 17504 88260 17508
rect 88196 17448 88246 17504
rect 88246 17448 88260 17504
rect 88196 17444 88260 17448
rect 93532 17504 93596 17508
rect 93532 17448 93582 17504
rect 93582 17448 93596 17504
rect 93532 17444 93596 17448
rect 122604 17444 122668 17508
rect 191052 17444 191116 17508
rect 253428 17444 253492 17508
rect 259500 17504 259564 17508
rect 259500 17448 259514 17504
rect 259514 17448 259564 17504
rect 259500 17444 259564 17448
rect 56916 17308 56980 17372
rect 65196 17308 65260 17372
rect 66300 17368 66364 17372
rect 66300 17312 66314 17368
rect 66314 17312 66364 17368
rect 66300 17308 66364 17312
rect 67588 17368 67652 17372
rect 67588 17312 67638 17368
rect 67638 17312 67652 17368
rect 67588 17308 67652 17312
rect 73292 17308 73356 17372
rect 98500 17308 98564 17372
rect 111012 17308 111076 17372
rect 248644 17308 248708 17372
rect 255820 17308 255884 17372
rect 256924 17308 256988 17372
rect 258396 17308 258460 17372
rect 35940 17172 36004 17236
rect 39620 17172 39684 17236
rect 61700 17172 61764 17236
rect 62804 17172 62868 17236
rect 63908 17172 63972 17236
rect 69796 17172 69860 17236
rect 70900 17172 70964 17236
rect 75684 17172 75748 17236
rect 192708 17172 192772 17236
rect 276060 17172 276124 17236
rect 283420 17172 283484 17236
rect 476068 17308 476132 17372
rect 472204 17172 472268 17236
rect 475700 17172 475764 17236
rect 58572 17036 58636 17100
rect 191788 17036 191852 17100
rect 251220 17096 251284 17100
rect 251220 17040 251234 17096
rect 251234 17040 251284 17096
rect 251220 17036 251284 17040
rect 414612 17036 414676 17100
rect 78260 16900 78324 16964
rect 465212 17036 465276 17100
rect 469628 17036 469692 17100
rect 478460 17036 478524 17100
rect 453620 16900 453684 16964
rect 478092 16900 478156 16964
rect 471284 16764 471348 16828
rect 416084 16628 416148 16692
rect 511028 16628 511092 16692
rect 357204 7652 357268 7716
rect 359964 7516 360028 7580
rect 419948 3708 420012 3772
rect 419764 3572 419828 3636
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 675244 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 675244 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 675244 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 675244 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 675244 49574 698058
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 675244 64454 676938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 675244 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 675244 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 675244 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 675244 85574 698058
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 675244 100454 676938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 675244 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 675244 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 675244 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 675244 121574 698058
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 675244 136454 676938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 675244 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 675244 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 675244 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 675244 157574 698058
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 150939 674932 151005 674933
rect 150939 674868 150940 674932
rect 151004 674868 151005 674932
rect 150939 674867 151005 674868
rect 150942 673470 151002 674867
rect 150840 673410 151002 673470
rect 150840 673202 150900 673410
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 20272 655174 20620 655206
rect 20272 654938 20328 655174
rect 20564 654938 20620 655174
rect 20272 654854 20620 654938
rect 20272 654618 20328 654854
rect 20564 654618 20620 654854
rect 20272 654586 20620 654618
rect 156000 655174 156348 655206
rect 156000 654938 156056 655174
rect 156292 654938 156348 655174
rect 156000 654854 156348 654938
rect 156000 654618 156056 654854
rect 156292 654618 156348 654854
rect 156000 654586 156348 654618
rect 20952 651454 21300 651486
rect 20952 651218 21008 651454
rect 21244 651218 21300 651454
rect 20952 651134 21300 651218
rect 20952 650898 21008 651134
rect 21244 650898 21300 651134
rect 20952 650866 21300 650898
rect 155320 651454 155668 651486
rect 155320 651218 155376 651454
rect 155612 651218 155668 651454
rect 155320 651134 155668 651218
rect 155320 650898 155376 651134
rect 155612 650898 155668 651134
rect 155320 650866 155668 650898
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 160674 630334 161294 665778
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 20272 619174 20620 619206
rect 20272 618938 20328 619174
rect 20564 618938 20620 619174
rect 20272 618854 20620 618938
rect 20272 618618 20328 618854
rect 20564 618618 20620 618854
rect 20272 618586 20620 618618
rect 156000 619174 156348 619206
rect 156000 618938 156056 619174
rect 156292 618938 156348 619174
rect 156000 618854 156348 618938
rect 156000 618618 156056 618854
rect 156292 618618 156348 618854
rect 156000 618586 156348 618618
rect 20952 615454 21300 615486
rect 20952 615218 21008 615454
rect 21244 615218 21300 615454
rect 20952 615134 21300 615218
rect 20952 614898 21008 615134
rect 21244 614898 21300 615134
rect 20952 614866 21300 614898
rect 155320 615454 155668 615486
rect 155320 615218 155376 615454
rect 155612 615218 155668 615454
rect 155320 615134 155668 615218
rect 155320 614898 155376 615134
rect 155612 614898 155668 615134
rect 155320 614866 155668 614898
rect 18643 598092 18709 598093
rect 18643 598028 18644 598092
rect 18708 598028 18709 598092
rect 18643 598027 18709 598028
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 17907 527236 17973 527237
rect 17907 527172 17908 527236
rect 17972 527172 17973 527236
rect 17907 527171 17973 527172
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 17910 521525 17970 527171
rect 17907 521524 17973 521525
rect 17907 521460 17908 521524
rect 17972 521460 17973 521524
rect 17907 521459 17973 521460
rect 18646 496093 18706 598027
rect 160674 594334 161294 629778
rect 160674 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 161294 594334
rect 160674 594014 161294 594098
rect 160674 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 161294 594014
rect 36056 589930 36116 590106
rect 37144 589930 37204 590106
rect 38232 589930 38292 590106
rect 35942 589870 36116 589930
rect 37046 589870 37204 589930
rect 38150 589870 38292 589930
rect 39592 589930 39652 590106
rect 40544 589930 40604 590106
rect 39592 589870 39682 589930
rect 35942 587757 36002 589870
rect 37046 587893 37106 589870
rect 37043 587892 37109 587893
rect 37043 587828 37044 587892
rect 37108 587828 37109 587892
rect 37043 587827 37109 587828
rect 35939 587756 36005 587757
rect 35939 587692 35940 587756
rect 36004 587692 36005 587756
rect 35939 587691 36005 587692
rect 38150 587621 38210 589870
rect 39622 587893 39682 589870
rect 40542 589870 40604 589930
rect 41768 589930 41828 590106
rect 43128 589930 43188 590106
rect 41768 589870 41890 589930
rect 39619 587892 39685 587893
rect 39619 587828 39620 587892
rect 39684 587828 39685 587892
rect 39619 587827 39685 587828
rect 19747 587620 19813 587621
rect 19747 587556 19748 587620
rect 19812 587556 19813 587620
rect 19747 587555 19813 587556
rect 38147 587620 38213 587621
rect 38147 587556 38148 587620
rect 38212 587556 38213 587620
rect 38147 587555 38213 587556
rect 19011 587348 19077 587349
rect 19011 587284 19012 587348
rect 19076 587284 19077 587348
rect 19011 587283 19077 587284
rect 18643 496092 18709 496093
rect 18643 496028 18644 496092
rect 18708 496028 18709 496092
rect 18643 496027 18709 496028
rect 19014 494733 19074 587283
rect 19011 494732 19077 494733
rect 19011 494668 19012 494732
rect 19076 494668 19077 494732
rect 19011 494667 19077 494668
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 18459 454340 18525 454341
rect 18459 454276 18460 454340
rect 18524 454276 18525 454340
rect 18459 454275 18525 454276
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 18462 96661 18522 454275
rect 19014 107405 19074 494667
rect 19750 491197 19810 587555
rect 40542 587485 40602 589870
rect 19931 587484 19997 587485
rect 19931 587420 19932 587484
rect 19996 587420 19997 587484
rect 19931 587419 19997 587420
rect 40539 587484 40605 587485
rect 40539 587420 40540 587484
rect 40604 587420 40605 587484
rect 40539 587419 40605 587420
rect 19934 497589 19994 587419
rect 41830 587349 41890 589870
rect 43118 589870 43188 589930
rect 44216 589930 44276 590106
rect 45440 589930 45500 590106
rect 44216 589870 44282 589930
rect 43118 587893 43178 589870
rect 44222 587893 44282 589870
rect 45326 589870 45500 589930
rect 46528 589930 46588 590106
rect 47616 589930 47676 590106
rect 48296 589930 48356 590106
rect 48704 589930 48764 590106
rect 46528 589870 46674 589930
rect 47616 589870 47778 589930
rect 45326 587893 45386 589870
rect 46614 587893 46674 589870
rect 47718 587893 47778 589870
rect 48270 589870 48356 589930
rect 48638 589870 48764 589930
rect 50064 589930 50124 590106
rect 50744 589930 50804 590106
rect 51288 589930 51348 590106
rect 52376 589930 52436 590106
rect 53464 589930 53524 590106
rect 50064 589870 50170 589930
rect 48270 587893 48330 589870
rect 43115 587892 43181 587893
rect 43115 587828 43116 587892
rect 43180 587828 43181 587892
rect 43115 587827 43181 587828
rect 44219 587892 44285 587893
rect 44219 587828 44220 587892
rect 44284 587828 44285 587892
rect 44219 587827 44285 587828
rect 45323 587892 45389 587893
rect 45323 587828 45324 587892
rect 45388 587828 45389 587892
rect 45323 587827 45389 587828
rect 46611 587892 46677 587893
rect 46611 587828 46612 587892
rect 46676 587828 46677 587892
rect 46611 587827 46677 587828
rect 47715 587892 47781 587893
rect 47715 587828 47716 587892
rect 47780 587828 47781 587892
rect 47715 587827 47781 587828
rect 48267 587892 48333 587893
rect 48267 587828 48268 587892
rect 48332 587828 48333 587892
rect 48267 587827 48333 587828
rect 48638 587757 48698 589870
rect 50110 587757 50170 589870
rect 50662 589870 50804 589930
rect 51214 589870 51348 589930
rect 52318 589870 52436 589930
rect 53422 589870 53524 589930
rect 53600 589930 53660 590106
rect 54552 589930 54612 590106
rect 55912 589930 55972 590106
rect 53600 589870 53666 589930
rect 50662 587893 50722 589870
rect 51214 587893 51274 589870
rect 52318 587893 52378 589870
rect 50659 587892 50725 587893
rect 50659 587828 50660 587892
rect 50724 587828 50725 587892
rect 50659 587827 50725 587828
rect 51211 587892 51277 587893
rect 51211 587828 51212 587892
rect 51276 587828 51277 587892
rect 51211 587827 51277 587828
rect 52315 587892 52381 587893
rect 52315 587828 52316 587892
rect 52380 587828 52381 587892
rect 52315 587827 52381 587828
rect 53422 587757 53482 589870
rect 53606 587893 53666 589870
rect 54526 589870 54612 589930
rect 55814 589870 55972 589930
rect 54526 587893 54586 589870
rect 55814 587893 55874 589870
rect 56048 589290 56108 590106
rect 57000 589930 57060 590106
rect 58088 589930 58148 590106
rect 58496 589930 58556 590106
rect 59448 589930 59508 590106
rect 60672 589930 60732 590106
rect 57000 589870 57162 589930
rect 58088 589870 58266 589930
rect 58496 589870 58634 589930
rect 59448 589870 59554 589930
rect 55998 589230 56108 589290
rect 55998 587893 56058 589230
rect 53603 587892 53669 587893
rect 53603 587828 53604 587892
rect 53668 587828 53669 587892
rect 53603 587827 53669 587828
rect 54523 587892 54589 587893
rect 54523 587828 54524 587892
rect 54588 587828 54589 587892
rect 54523 587827 54589 587828
rect 55811 587892 55877 587893
rect 55811 587828 55812 587892
rect 55876 587828 55877 587892
rect 55811 587827 55877 587828
rect 55995 587892 56061 587893
rect 55995 587828 55996 587892
rect 56060 587828 56061 587892
rect 55995 587827 56061 587828
rect 48635 587756 48701 587757
rect 48635 587692 48636 587756
rect 48700 587692 48701 587756
rect 48635 587691 48701 587692
rect 50107 587756 50173 587757
rect 50107 587692 50108 587756
rect 50172 587692 50173 587756
rect 50107 587691 50173 587692
rect 53419 587756 53485 587757
rect 53419 587692 53420 587756
rect 53484 587692 53485 587756
rect 53419 587691 53485 587692
rect 57102 587485 57162 589870
rect 58206 587621 58266 589870
rect 58574 587893 58634 589870
rect 58571 587892 58637 587893
rect 58571 587828 58572 587892
rect 58636 587828 58637 587892
rect 58571 587827 58637 587828
rect 59494 587757 59554 589870
rect 60598 589870 60732 589930
rect 61080 589930 61140 590106
rect 61760 589930 61820 590106
rect 62848 589930 62908 590106
rect 61080 589870 61210 589930
rect 60598 587893 60658 589870
rect 60595 587892 60661 587893
rect 60595 587828 60596 587892
rect 60660 587828 60661 587892
rect 60595 587827 60661 587828
rect 59491 587756 59557 587757
rect 59491 587692 59492 587756
rect 59556 587692 59557 587756
rect 59491 587691 59557 587692
rect 58203 587620 58269 587621
rect 58203 587556 58204 587620
rect 58268 587556 58269 587620
rect 58203 587555 58269 587556
rect 57099 587484 57165 587485
rect 57099 587420 57100 587484
rect 57164 587420 57165 587484
rect 57099 587419 57165 587420
rect 41827 587348 41893 587349
rect 41827 587284 41828 587348
rect 41892 587284 41893 587348
rect 41827 587283 41893 587284
rect 58206 587213 58266 587555
rect 61150 587349 61210 589870
rect 61702 589870 61820 589930
rect 62806 589870 62908 589930
rect 63528 589930 63588 590106
rect 63936 589930 63996 590106
rect 65296 589930 65356 590106
rect 65976 589930 66036 590106
rect 66384 589930 66444 590106
rect 67608 589930 67668 590106
rect 63528 589870 63602 589930
rect 61702 587893 61762 589870
rect 62806 587893 62866 589870
rect 61699 587892 61765 587893
rect 61699 587828 61700 587892
rect 61764 587828 61765 587892
rect 61699 587827 61765 587828
rect 62803 587892 62869 587893
rect 62803 587828 62804 587892
rect 62868 587828 62869 587892
rect 62803 587827 62869 587828
rect 63542 587349 63602 589870
rect 63910 589870 63996 589930
rect 65198 589870 65356 589930
rect 65934 589870 66036 589930
rect 66302 589870 66444 589930
rect 67590 589870 67668 589930
rect 68288 589930 68348 590106
rect 68696 589930 68756 590106
rect 68288 589870 68386 589930
rect 63910 587893 63970 589870
rect 65198 587893 65258 589870
rect 63907 587892 63973 587893
rect 63907 587828 63908 587892
rect 63972 587828 63973 587892
rect 63907 587827 63973 587828
rect 65195 587892 65261 587893
rect 65195 587828 65196 587892
rect 65260 587828 65261 587892
rect 65195 587827 65261 587828
rect 65934 587485 65994 589870
rect 66302 587893 66362 589870
rect 67590 587893 67650 589870
rect 66299 587892 66365 587893
rect 66299 587828 66300 587892
rect 66364 587828 66365 587892
rect 66299 587827 66365 587828
rect 67587 587892 67653 587893
rect 67587 587828 67588 587892
rect 67652 587828 67653 587892
rect 67587 587827 67653 587828
rect 68326 587485 68386 589870
rect 68694 589870 68756 589930
rect 69784 589930 69844 590106
rect 71008 589930 71068 590106
rect 69784 589870 69858 589930
rect 68694 587893 68754 589870
rect 69798 587893 69858 589870
rect 70902 589870 71068 589930
rect 71144 589930 71204 590106
rect 72232 589930 72292 590106
rect 73320 589930 73380 590106
rect 71144 589870 71330 589930
rect 68691 587892 68757 587893
rect 68691 587828 68692 587892
rect 68756 587828 68757 587892
rect 68691 587827 68757 587828
rect 69795 587892 69861 587893
rect 69795 587828 69796 587892
rect 69860 587828 69861 587892
rect 69795 587827 69861 587828
rect 65931 587484 65997 587485
rect 65931 587420 65932 587484
rect 65996 587420 65997 587484
rect 65931 587419 65997 587420
rect 68323 587484 68389 587485
rect 68323 587420 68324 587484
rect 68388 587420 68389 587484
rect 68323 587419 68389 587420
rect 61147 587348 61213 587349
rect 61147 587284 61148 587348
rect 61212 587284 61213 587348
rect 61147 587283 61213 587284
rect 63539 587348 63605 587349
rect 63539 587284 63540 587348
rect 63604 587284 63605 587348
rect 63539 587283 63605 587284
rect 70902 587213 70962 589870
rect 71270 587893 71330 589870
rect 72190 589870 72292 589930
rect 73294 589870 73380 589930
rect 73592 589930 73652 590106
rect 74408 589930 74468 590106
rect 75768 589930 75828 590106
rect 73592 589870 73722 589930
rect 72190 587893 72250 589870
rect 73294 587893 73354 589870
rect 73662 587893 73722 589870
rect 74398 589870 74468 589930
rect 75686 589870 75828 589930
rect 74398 587893 74458 589870
rect 71267 587892 71333 587893
rect 71267 587828 71268 587892
rect 71332 587828 71333 587892
rect 71267 587827 71333 587828
rect 72187 587892 72253 587893
rect 72187 587828 72188 587892
rect 72252 587828 72253 587892
rect 72187 587827 72253 587828
rect 73291 587892 73357 587893
rect 73291 587828 73292 587892
rect 73356 587828 73357 587892
rect 73291 587827 73357 587828
rect 73659 587892 73725 587893
rect 73659 587828 73660 587892
rect 73724 587828 73725 587892
rect 73659 587827 73725 587828
rect 74395 587892 74461 587893
rect 74395 587828 74396 587892
rect 74460 587828 74461 587892
rect 74395 587827 74461 587828
rect 75686 587621 75746 589870
rect 76040 589658 76100 590106
rect 76992 589658 77052 590106
rect 78080 589658 78140 590106
rect 78488 589658 78548 590106
rect 76040 589598 76114 589658
rect 76054 587893 76114 589598
rect 76974 589598 77052 589658
rect 78078 589598 78140 589658
rect 78446 589598 78548 589658
rect 79168 589658 79228 590106
rect 80936 589930 80996 590106
rect 83520 589930 83580 590106
rect 85968 589930 86028 590106
rect 88280 589930 88340 590106
rect 91000 589930 91060 590106
rect 80936 589870 81082 589930
rect 83520 589870 83658 589930
rect 85968 589870 86050 589930
rect 79168 589598 79242 589658
rect 76051 587892 76117 587893
rect 76051 587828 76052 587892
rect 76116 587828 76117 587892
rect 76051 587827 76117 587828
rect 75683 587620 75749 587621
rect 75683 587556 75684 587620
rect 75748 587556 75749 587620
rect 75683 587555 75749 587556
rect 76974 587485 77034 589598
rect 78078 587893 78138 589598
rect 78446 587893 78506 589598
rect 79182 587893 79242 589598
rect 81022 587893 81082 589870
rect 83598 587893 83658 589870
rect 78075 587892 78141 587893
rect 78075 587828 78076 587892
rect 78140 587828 78141 587892
rect 78075 587827 78141 587828
rect 78443 587892 78509 587893
rect 78443 587828 78444 587892
rect 78508 587828 78509 587892
rect 78443 587827 78509 587828
rect 79179 587892 79245 587893
rect 79179 587828 79180 587892
rect 79244 587828 79245 587892
rect 79179 587827 79245 587828
rect 81019 587892 81085 587893
rect 81019 587828 81020 587892
rect 81084 587828 81085 587892
rect 81019 587827 81085 587828
rect 83595 587892 83661 587893
rect 83595 587828 83596 587892
rect 83660 587828 83661 587892
rect 83595 587827 83661 587828
rect 76971 587484 77037 587485
rect 76971 587420 76972 587484
rect 77036 587420 77037 587484
rect 76971 587419 77037 587420
rect 85990 587349 86050 589870
rect 88198 589870 88340 589930
rect 90958 589870 91060 589930
rect 93448 589930 93508 590106
rect 95896 589930 95956 590106
rect 98480 589930 98540 590106
rect 100928 589930 100988 590106
rect 103512 589930 103572 590106
rect 105960 589930 106020 590106
rect 108544 589930 108604 590106
rect 93448 589870 93594 589930
rect 95896 589870 95986 589930
rect 98480 589870 98562 589930
rect 88198 587893 88258 589870
rect 90958 587893 91018 589870
rect 93534 587893 93594 589870
rect 95926 587893 95986 589870
rect 98502 587893 98562 589870
rect 100894 589870 100988 589930
rect 103286 589870 103572 589930
rect 105862 589870 106020 589930
rect 108438 589870 108604 589930
rect 110992 589930 111052 590106
rect 113440 589930 113500 590106
rect 115888 589930 115948 590106
rect 118472 589930 118532 590106
rect 110992 589870 111074 589930
rect 100894 587893 100954 589870
rect 88195 587892 88261 587893
rect 88195 587828 88196 587892
rect 88260 587828 88261 587892
rect 88195 587827 88261 587828
rect 90955 587892 91021 587893
rect 90955 587828 90956 587892
rect 91020 587828 91021 587892
rect 90955 587827 91021 587828
rect 93531 587892 93597 587893
rect 93531 587828 93532 587892
rect 93596 587828 93597 587892
rect 93531 587827 93597 587828
rect 95923 587892 95989 587893
rect 95923 587828 95924 587892
rect 95988 587828 95989 587892
rect 95923 587827 95989 587828
rect 98499 587892 98565 587893
rect 98499 587828 98500 587892
rect 98564 587828 98565 587892
rect 98499 587827 98565 587828
rect 100891 587892 100957 587893
rect 100891 587828 100892 587892
rect 100956 587828 100957 587892
rect 103286 587890 103346 589870
rect 105862 587893 105922 589870
rect 108438 587893 108498 589870
rect 111014 587893 111074 589870
rect 113406 589870 113500 589930
rect 115798 589870 115948 589930
rect 118374 589870 118532 589930
rect 120920 589930 120980 590106
rect 123368 589930 123428 590106
rect 125952 589930 126012 590106
rect 120920 589870 121010 589930
rect 113406 587893 113466 589870
rect 115798 587893 115858 589870
rect 118374 587893 118434 589870
rect 120950 587893 121010 589870
rect 123342 589870 123428 589930
rect 125918 589870 126012 589930
rect 123342 589290 123402 589870
rect 122606 589230 123402 589290
rect 103467 587892 103533 587893
rect 103467 587890 103468 587892
rect 103286 587830 103468 587890
rect 100891 587827 100957 587828
rect 103467 587828 103468 587830
rect 103532 587828 103533 587892
rect 103467 587827 103533 587828
rect 105859 587892 105925 587893
rect 105859 587828 105860 587892
rect 105924 587828 105925 587892
rect 105859 587827 105925 587828
rect 108435 587892 108501 587893
rect 108435 587828 108436 587892
rect 108500 587828 108501 587892
rect 108435 587827 108501 587828
rect 111011 587892 111077 587893
rect 111011 587828 111012 587892
rect 111076 587828 111077 587892
rect 111011 587827 111077 587828
rect 113403 587892 113469 587893
rect 113403 587828 113404 587892
rect 113468 587828 113469 587892
rect 113403 587827 113469 587828
rect 115795 587892 115861 587893
rect 115795 587828 115796 587892
rect 115860 587828 115861 587892
rect 115795 587827 115861 587828
rect 118371 587892 118437 587893
rect 118371 587828 118372 587892
rect 118436 587828 118437 587892
rect 118371 587827 118437 587828
rect 120947 587892 121013 587893
rect 120947 587828 120948 587892
rect 121012 587828 121013 587892
rect 120947 587827 121013 587828
rect 85987 587348 86053 587349
rect 85987 587284 85988 587348
rect 86052 587284 86053 587348
rect 85987 587283 86053 587284
rect 58203 587212 58269 587213
rect 58203 587148 58204 587212
rect 58268 587148 58269 587212
rect 58203 587147 58269 587148
rect 70899 587212 70965 587213
rect 70899 587148 70900 587212
rect 70964 587148 70965 587212
rect 122606 587210 122666 589230
rect 125918 587893 125978 589870
rect 125915 587892 125981 587893
rect 125915 587828 125916 587892
rect 125980 587828 125981 587892
rect 125915 587827 125981 587828
rect 122606 587150 122850 587210
rect 70899 587147 70965 587148
rect 122790 587077 122850 587150
rect 122787 587076 122853 587077
rect 122787 587012 122788 587076
rect 122852 587012 122853 587076
rect 122787 587011 122853 587012
rect 150755 585308 150821 585309
rect 150755 585244 150756 585308
rect 150820 585244 150821 585308
rect 150755 585243 150821 585244
rect 150758 583810 150818 585243
rect 150758 583750 150900 583810
rect 150840 583202 150900 583750
rect 20272 582929 20620 583036
rect 20272 582693 20328 582929
rect 20564 582693 20620 582929
rect 20272 582586 20620 582693
rect 156000 582929 156348 583036
rect 156000 582693 156056 582929
rect 156292 582693 156348 582929
rect 156000 582586 156348 582693
rect 20952 579454 21300 579486
rect 20952 579218 21008 579454
rect 21244 579218 21300 579454
rect 20952 579134 21300 579218
rect 20952 578898 21008 579134
rect 21244 578898 21300 579134
rect 20952 578866 21300 578898
rect 155320 579454 155668 579486
rect 155320 579218 155376 579454
rect 155612 579218 155668 579454
rect 155320 579134 155668 579218
rect 155320 578898 155376 579134
rect 155612 578898 155668 579134
rect 155320 578866 155668 578898
rect 160674 558334 161294 593778
rect 160674 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 161294 558334
rect 160674 558014 161294 558098
rect 160674 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 161294 558014
rect 20272 547174 20620 547206
rect 20272 546938 20328 547174
rect 20564 546938 20620 547174
rect 20272 546854 20620 546938
rect 20272 546618 20328 546854
rect 20564 546618 20620 546854
rect 20272 546586 20620 546618
rect 156000 547174 156348 547206
rect 156000 546938 156056 547174
rect 156292 546938 156348 547174
rect 156000 546854 156348 546938
rect 156000 546618 156056 546854
rect 156292 546618 156348 546854
rect 156000 546586 156348 546618
rect 20952 543454 21300 543486
rect 20952 543218 21008 543454
rect 21244 543218 21300 543454
rect 20952 543134 21300 543218
rect 20952 542898 21008 543134
rect 21244 542898 21300 543134
rect 20952 542866 21300 542898
rect 155320 543454 155668 543486
rect 155320 543218 155376 543454
rect 155612 543218 155668 543454
rect 155320 543134 155668 543218
rect 155320 542898 155376 543134
rect 155612 542898 155668 543134
rect 155320 542866 155668 542898
rect 160674 522334 161294 557778
rect 160674 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 161294 522334
rect 160674 522014 161294 522098
rect 160674 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 161294 522014
rect 20272 511174 20620 511206
rect 20272 510938 20328 511174
rect 20564 510938 20620 511174
rect 20272 510854 20620 510938
rect 20272 510618 20328 510854
rect 20564 510618 20620 510854
rect 20272 510586 20620 510618
rect 156000 511174 156348 511206
rect 156000 510938 156056 511174
rect 156292 510938 156348 511174
rect 156000 510854 156348 510938
rect 156000 510618 156056 510854
rect 156292 510618 156348 510854
rect 156000 510586 156348 510618
rect 20952 507454 21300 507486
rect 20952 507218 21008 507454
rect 21244 507218 21300 507454
rect 20952 507134 21300 507218
rect 20952 506898 21008 507134
rect 21244 506898 21300 507134
rect 20952 506866 21300 506898
rect 155320 507454 155668 507486
rect 155320 507218 155376 507454
rect 155612 507218 155668 507454
rect 155320 507134 155668 507218
rect 155320 506898 155376 507134
rect 155612 506898 155668 507134
rect 155320 506866 155668 506898
rect 36056 499590 36116 500106
rect 37144 499590 37204 500106
rect 38232 499590 38292 500106
rect 36056 499530 36186 499590
rect 37144 499530 37290 499590
rect 19931 497588 19997 497589
rect 19931 497524 19932 497588
rect 19996 497524 19997 497588
rect 19931 497523 19997 497524
rect 19747 491196 19813 491197
rect 19747 491132 19748 491196
rect 19812 491132 19813 491196
rect 19747 491131 19813 491132
rect 19195 456924 19261 456925
rect 19195 456860 19196 456924
rect 19260 456860 19261 456924
rect 19195 456859 19261 456860
rect 19011 107404 19077 107405
rect 19011 107340 19012 107404
rect 19076 107340 19077 107404
rect 19011 107339 19077 107340
rect 18459 96660 18525 96661
rect 18459 96596 18460 96660
rect 18524 96596 18525 96660
rect 18459 96595 18525 96596
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 19014 17781 19074 107339
rect 19198 28117 19258 456859
rect 19934 107541 19994 497523
rect 20394 490054 21014 498064
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 195244 21014 201498
rect 24114 493774 24734 498064
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 24114 195244 24734 205218
rect 27834 497494 28454 498064
rect 36126 497861 36186 499530
rect 37230 497861 37290 499530
rect 38150 499530 38292 499590
rect 39592 499590 39652 500106
rect 40544 499590 40604 500106
rect 39592 499530 39682 499590
rect 38150 498133 38210 499530
rect 38147 498132 38213 498133
rect 38147 498068 38148 498132
rect 38212 498068 38213 498132
rect 38147 498067 38213 498068
rect 36123 497860 36189 497861
rect 36123 497796 36124 497860
rect 36188 497796 36189 497860
rect 36123 497795 36189 497796
rect 37227 497860 37293 497861
rect 37227 497796 37228 497860
rect 37292 497796 37293 497860
rect 37227 497795 37293 497796
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 27834 195244 28454 208938
rect 37794 471454 38414 497940
rect 39622 497045 39682 499530
rect 40542 499530 40604 499590
rect 41768 499590 41828 500106
rect 43128 499590 43188 500106
rect 41768 499530 41890 499590
rect 39619 497044 39685 497045
rect 39619 496980 39620 497044
rect 39684 496980 39685 497044
rect 39619 496979 39685 496980
rect 40542 496909 40602 499530
rect 41830 498133 41890 499530
rect 43118 499530 43188 499590
rect 44216 499590 44276 500106
rect 45440 499629 45500 500106
rect 45437 499628 45503 499629
rect 44216 499530 44282 499590
rect 45437 499564 45438 499628
rect 45502 499564 45503 499628
rect 45437 499563 45503 499564
rect 46528 499590 46588 500106
rect 47616 499590 47676 500106
rect 48296 499590 48356 500106
rect 48704 499590 48764 500106
rect 46528 499530 46674 499590
rect 43118 498133 43178 499530
rect 41827 498132 41893 498133
rect 41827 498068 41828 498132
rect 41892 498068 41893 498132
rect 41827 498067 41893 498068
rect 43115 498132 43181 498133
rect 43115 498068 43116 498132
rect 43180 498068 43181 498132
rect 43115 498067 43181 498068
rect 44222 497997 44282 499530
rect 46614 498133 46674 499530
rect 47534 499530 47676 499590
rect 48270 499530 48356 499590
rect 48638 499530 48764 499590
rect 50064 499590 50124 500106
rect 50744 499590 50804 500106
rect 51288 499590 51348 500106
rect 52376 499590 52436 500106
rect 53464 499590 53524 500106
rect 50064 499530 50170 499590
rect 50744 499530 50906 499590
rect 51288 499530 51458 499590
rect 47534 498133 47594 499530
rect 46611 498132 46677 498133
rect 46611 498068 46612 498132
rect 46676 498068 46677 498132
rect 46611 498067 46677 498068
rect 47531 498132 47597 498133
rect 47531 498068 47532 498132
rect 47596 498068 47597 498132
rect 47531 498067 47597 498068
rect 44219 497996 44285 497997
rect 40539 496908 40605 496909
rect 40539 496844 40540 496908
rect 40604 496844 40605 496908
rect 40539 496843 40605 496844
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 195244 38414 218898
rect 41514 475174 42134 497940
rect 44219 497932 44220 497996
rect 44284 497932 44285 497996
rect 44219 497931 44285 497932
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 195244 42134 222618
rect 45234 478894 45854 497940
rect 48270 496909 48330 499530
rect 48638 498133 48698 499530
rect 48635 498132 48701 498133
rect 48635 498068 48636 498132
rect 48700 498068 48701 498132
rect 48635 498067 48701 498068
rect 48267 496908 48333 496909
rect 48267 496844 48268 496908
rect 48332 496844 48333 496908
rect 48267 496843 48333 496844
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 195244 45854 226338
rect 48954 482614 49574 498064
rect 50110 497861 50170 499530
rect 50107 497860 50173 497861
rect 50107 497796 50108 497860
rect 50172 497796 50173 497860
rect 50107 497795 50173 497796
rect 50846 496909 50906 499530
rect 51398 498133 51458 499530
rect 52318 499530 52436 499590
rect 53422 499530 53524 499590
rect 53600 499590 53660 500106
rect 54552 499590 54612 500106
rect 55912 499590 55972 500106
rect 53600 499530 53666 499590
rect 52318 498133 52378 499530
rect 53422 498133 53482 499530
rect 51395 498132 51461 498133
rect 51395 498068 51396 498132
rect 51460 498068 51461 498132
rect 51395 498067 51461 498068
rect 52315 498132 52381 498133
rect 52315 498068 52316 498132
rect 52380 498068 52381 498132
rect 52315 498067 52381 498068
rect 53419 498132 53485 498133
rect 53419 498068 53420 498132
rect 53484 498068 53485 498132
rect 53419 498067 53485 498068
rect 50843 496908 50909 496909
rect 50843 496844 50844 496908
rect 50908 496844 50909 496908
rect 50843 496843 50909 496844
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 195244 49574 230058
rect 52674 486334 53294 498064
rect 53606 496909 53666 499530
rect 54526 499530 54612 499590
rect 55814 499530 55972 499590
rect 56048 499590 56108 500106
rect 57000 499590 57060 500106
rect 58088 499590 58148 500106
rect 58496 499590 58556 500106
rect 59448 499590 59508 500106
rect 60672 499590 60732 500106
rect 56048 499530 56242 499590
rect 57000 499530 57162 499590
rect 58088 499530 58266 499590
rect 58496 499530 58634 499590
rect 59448 499530 59554 499590
rect 54526 498133 54586 499530
rect 55814 498133 55874 499530
rect 54523 498132 54589 498133
rect 54523 498068 54524 498132
rect 54588 498068 54589 498132
rect 54523 498067 54589 498068
rect 55811 498132 55877 498133
rect 55811 498068 55812 498132
rect 55876 498068 55877 498132
rect 55811 498067 55877 498068
rect 56182 496909 56242 499530
rect 53603 496908 53669 496909
rect 53603 496844 53604 496908
rect 53668 496844 53669 496908
rect 53603 496843 53669 496844
rect 56179 496908 56245 496909
rect 56179 496844 56180 496908
rect 56244 496844 56245 496908
rect 56179 496843 56245 496844
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52674 414334 53294 449778
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52674 378334 53294 413778
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 52674 342334 53294 377778
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52674 306334 53294 341778
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52674 270334 53294 305778
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52674 234334 53294 269778
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52674 198334 53294 233778
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52674 195244 53294 197778
rect 56394 490054 57014 497940
rect 57102 497861 57162 499530
rect 58206 497997 58266 499530
rect 58203 497996 58269 497997
rect 58203 497932 58204 497996
rect 58268 497932 58269 497996
rect 58203 497931 58269 497932
rect 57099 497860 57165 497861
rect 57099 497796 57100 497860
rect 57164 497796 57165 497860
rect 57099 497795 57165 497796
rect 58574 496909 58634 499530
rect 59494 498133 59554 499530
rect 60598 499530 60732 499590
rect 61080 499590 61140 500106
rect 61760 499590 61820 500106
rect 62848 499590 62908 500106
rect 61080 499530 61210 499590
rect 60598 498133 60658 499530
rect 59491 498132 59557 498133
rect 59491 498068 59492 498132
rect 59556 498068 59557 498132
rect 59491 498067 59557 498068
rect 60595 498132 60661 498133
rect 60595 498068 60596 498132
rect 60660 498068 60661 498132
rect 60595 498067 60661 498068
rect 58571 496908 58637 496909
rect 58571 496844 58572 496908
rect 58636 496844 58637 496908
rect 58571 496843 58637 496844
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 56394 454054 57014 489498
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 56394 418054 57014 453498
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 56394 382054 57014 417498
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 56394 346054 57014 381498
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 56394 310054 57014 345498
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 56394 274054 57014 309498
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 56394 238054 57014 273498
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 56394 202054 57014 237498
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 195244 57014 201498
rect 60114 493774 60734 497940
rect 61150 496909 61210 499530
rect 61702 499530 61820 499590
rect 62806 499530 62908 499590
rect 63528 499590 63588 500106
rect 63936 499590 63996 500106
rect 63528 499530 63602 499590
rect 61702 497045 61762 499530
rect 61699 497044 61765 497045
rect 61699 496980 61700 497044
rect 61764 496980 61765 497044
rect 61699 496979 61765 496980
rect 62806 496909 62866 499530
rect 63542 498133 63602 499530
rect 63910 499530 63996 499590
rect 65296 499590 65356 500106
rect 65976 499590 66036 500106
rect 66384 499590 66444 500106
rect 67608 499590 67668 500106
rect 65296 499530 65442 499590
rect 63910 498133 63970 499530
rect 63539 498132 63605 498133
rect 63539 498068 63540 498132
rect 63604 498068 63605 498132
rect 63539 498067 63605 498068
rect 63907 498132 63973 498133
rect 63907 498068 63908 498132
rect 63972 498068 63973 498132
rect 63907 498067 63973 498068
rect 63834 497494 64454 497940
rect 63834 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 64454 497494
rect 63834 497174 64454 497258
rect 63834 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 64454 497174
rect 61147 496908 61213 496909
rect 61147 496844 61148 496908
rect 61212 496844 61213 496908
rect 61147 496843 61213 496844
rect 62803 496908 62869 496909
rect 62803 496844 62804 496908
rect 62868 496844 62869 496908
rect 62803 496843 62869 496844
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 60114 421774 60734 457218
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 60114 385774 60734 421218
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 60114 349774 60734 385218
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 313774 60734 349218
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 60114 277774 60734 313218
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 60114 241774 60734 277218
rect 60114 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 60734 241774
rect 60114 241454 60734 241538
rect 60114 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 60734 241454
rect 60114 205774 60734 241218
rect 60114 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 60734 205774
rect 60114 205454 60734 205538
rect 60114 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 60734 205454
rect 60114 195244 60734 205218
rect 63834 461494 64454 496938
rect 65382 496909 65442 499530
rect 65934 499530 66036 499590
rect 66302 499530 66444 499590
rect 67590 499530 67668 499590
rect 68288 499590 68348 500106
rect 68696 499590 68756 500106
rect 68288 499530 68386 499590
rect 65934 496909 65994 499530
rect 66302 497045 66362 499530
rect 67590 498133 67650 499530
rect 67587 498132 67653 498133
rect 67587 498068 67588 498132
rect 67652 498068 67653 498132
rect 67587 498067 67653 498068
rect 66299 497044 66365 497045
rect 66299 496980 66300 497044
rect 66364 496980 66365 497044
rect 66299 496979 66365 496980
rect 68326 496909 68386 499530
rect 68694 499530 68756 499590
rect 69784 499590 69844 500106
rect 71008 499590 71068 500106
rect 69784 499530 69858 499590
rect 68694 497181 68754 499530
rect 68691 497180 68757 497181
rect 68691 497116 68692 497180
rect 68756 497116 68757 497180
rect 68691 497115 68757 497116
rect 69798 496909 69858 499530
rect 70902 499530 71068 499590
rect 71144 499590 71204 500106
rect 72232 499590 72292 500106
rect 73320 499590 73380 500106
rect 71144 499530 71330 499590
rect 70902 496909 70962 499530
rect 71270 498133 71330 499530
rect 72190 499530 72292 499590
rect 73294 499530 73380 499590
rect 73592 499590 73652 500106
rect 74408 499590 74468 500106
rect 75768 499590 75828 500106
rect 73592 499530 73722 499590
rect 72190 498133 72250 499530
rect 71267 498132 71333 498133
rect 71267 498068 71268 498132
rect 71332 498068 71333 498132
rect 71267 498067 71333 498068
rect 72187 498132 72253 498133
rect 72187 498068 72188 498132
rect 72252 498068 72253 498132
rect 72187 498067 72253 498068
rect 73294 497725 73354 499530
rect 73662 498133 73722 499530
rect 74398 499530 74468 499590
rect 75686 499530 75828 499590
rect 76040 499590 76100 500106
rect 76992 499590 77052 500106
rect 78080 499590 78140 500106
rect 78488 499590 78548 500106
rect 76040 499530 76114 499590
rect 74398 498133 74458 499530
rect 73659 498132 73725 498133
rect 73659 498068 73660 498132
rect 73724 498068 73725 498132
rect 73659 498067 73725 498068
rect 74395 498132 74461 498133
rect 74395 498068 74396 498132
rect 74460 498068 74461 498132
rect 74395 498067 74461 498068
rect 73291 497724 73357 497725
rect 73291 497660 73292 497724
rect 73356 497660 73357 497724
rect 73291 497659 73357 497660
rect 73294 496909 73354 497659
rect 65379 496908 65445 496909
rect 65379 496844 65380 496908
rect 65444 496844 65445 496908
rect 65379 496843 65445 496844
rect 65931 496908 65997 496909
rect 65931 496844 65932 496908
rect 65996 496844 65997 496908
rect 65931 496843 65997 496844
rect 68323 496908 68389 496909
rect 68323 496844 68324 496908
rect 68388 496844 68389 496908
rect 68323 496843 68389 496844
rect 69795 496908 69861 496909
rect 69795 496844 69796 496908
rect 69860 496844 69861 496908
rect 69795 496843 69861 496844
rect 70899 496908 70965 496909
rect 70899 496844 70900 496908
rect 70964 496844 70965 496908
rect 70899 496843 70965 496844
rect 73291 496908 73357 496909
rect 73291 496844 73292 496908
rect 73356 496844 73357 496908
rect 73291 496843 73357 496844
rect 63834 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 64454 461494
rect 63834 461174 64454 461258
rect 63834 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 64454 461174
rect 63834 425494 64454 460938
rect 63834 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 64454 425494
rect 63834 425174 64454 425258
rect 63834 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 64454 425174
rect 63834 389494 64454 424938
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 63834 353494 64454 388938
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63834 317494 64454 352938
rect 63834 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 64454 317494
rect 63834 317174 64454 317258
rect 63834 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 64454 317174
rect 63834 281494 64454 316938
rect 63834 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 64454 281494
rect 63834 281174 64454 281258
rect 63834 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 64454 281174
rect 63834 245494 64454 280938
rect 63834 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 64454 245494
rect 63834 245174 64454 245258
rect 63834 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 64454 245174
rect 63834 209494 64454 244938
rect 63834 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 64454 209494
rect 63834 209174 64454 209258
rect 63834 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 64454 209174
rect 63834 195244 64454 208938
rect 73794 471454 74414 497940
rect 75686 497861 75746 499530
rect 75683 497860 75749 497861
rect 75683 497796 75684 497860
rect 75748 497796 75749 497860
rect 75683 497795 75749 497796
rect 76054 496909 76114 499530
rect 76974 499530 77052 499590
rect 78078 499530 78140 499590
rect 78446 499530 78548 499590
rect 79168 499590 79228 500106
rect 80936 499590 80996 500106
rect 83520 499590 83580 500106
rect 85968 499590 86028 500106
rect 88280 499590 88340 500106
rect 91000 499590 91060 500106
rect 79168 499530 79242 499590
rect 80936 499530 81082 499590
rect 83520 499530 83658 499590
rect 85968 499530 86050 499590
rect 76974 497997 77034 499530
rect 78078 498133 78138 499530
rect 78075 498132 78141 498133
rect 78075 498068 78076 498132
rect 78140 498068 78141 498132
rect 78075 498067 78141 498068
rect 76971 497996 77037 497997
rect 76971 497932 76972 497996
rect 77036 497932 77037 497996
rect 76971 497931 77037 497932
rect 76051 496908 76117 496909
rect 76051 496844 76052 496908
rect 76116 496844 76117 496908
rect 76051 496843 76117 496844
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 195244 74414 218898
rect 77514 475174 78134 497940
rect 78446 496909 78506 499530
rect 79182 496909 79242 499530
rect 81022 496909 81082 499530
rect 78443 496908 78509 496909
rect 78443 496844 78444 496908
rect 78508 496844 78509 496908
rect 78443 496843 78509 496844
rect 79179 496908 79245 496909
rect 79179 496844 79180 496908
rect 79244 496844 79245 496908
rect 79179 496843 79245 496844
rect 81019 496908 81085 496909
rect 81019 496844 81020 496908
rect 81084 496844 81085 496908
rect 81019 496843 81085 496844
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 195244 78134 222618
rect 81234 478894 81854 498064
rect 83598 496909 83658 499530
rect 83595 496908 83661 496909
rect 83595 496844 83596 496908
rect 83660 496844 83661 496908
rect 83595 496843 83661 496844
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 195244 81854 226338
rect 84954 482614 85574 498064
rect 85990 496909 86050 499530
rect 88198 499530 88340 499590
rect 90958 499530 91060 499590
rect 93448 499590 93508 500106
rect 95896 499590 95956 500106
rect 98480 499590 98540 500106
rect 100928 499590 100988 500106
rect 93448 499530 93594 499590
rect 95896 499530 95986 499590
rect 98480 499530 98562 499590
rect 88198 496909 88258 499530
rect 85987 496908 86053 496909
rect 85987 496844 85988 496908
rect 86052 496844 86053 496908
rect 85987 496843 86053 496844
rect 88195 496908 88261 496909
rect 88195 496844 88196 496908
rect 88260 496844 88261 496908
rect 88195 496843 88261 496844
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 195244 85574 230058
rect 88674 486334 89294 498064
rect 90958 496909 91018 499530
rect 90955 496908 91021 496909
rect 90955 496844 90956 496908
rect 91020 496844 91021 496908
rect 90955 496843 91021 496844
rect 88674 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 89294 486334
rect 88674 486014 89294 486098
rect 88674 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 89294 486014
rect 88674 450334 89294 485778
rect 88674 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 89294 450334
rect 88674 450014 89294 450098
rect 88674 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 89294 450014
rect 88674 414334 89294 449778
rect 88674 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 89294 414334
rect 88674 414014 89294 414098
rect 88674 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 89294 414014
rect 88674 378334 89294 413778
rect 88674 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 89294 378334
rect 88674 378014 89294 378098
rect 88674 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 89294 378014
rect 88674 342334 89294 377778
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 88674 306334 89294 341778
rect 88674 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 89294 306334
rect 88674 306014 89294 306098
rect 88674 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 89294 306014
rect 88674 270334 89294 305778
rect 88674 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 89294 270334
rect 88674 270014 89294 270098
rect 88674 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 89294 270014
rect 88674 234334 89294 269778
rect 88674 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 89294 234334
rect 88674 234014 89294 234098
rect 88674 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 89294 234014
rect 88674 198334 89294 233778
rect 88674 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 89294 198334
rect 88674 198014 89294 198098
rect 88674 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 89294 198014
rect 88674 195244 89294 197778
rect 92394 490054 93014 498064
rect 93534 496909 93594 499530
rect 95926 496909 95986 499530
rect 93531 496908 93597 496909
rect 93531 496844 93532 496908
rect 93596 496844 93597 496908
rect 93531 496843 93597 496844
rect 95923 496908 95989 496909
rect 95923 496844 95924 496908
rect 95988 496844 95989 496908
rect 95923 496843 95989 496844
rect 92394 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 93014 490054
rect 92394 489734 93014 489818
rect 92394 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 93014 489734
rect 92394 454054 93014 489498
rect 92394 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 93014 454054
rect 92394 453734 93014 453818
rect 92394 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 93014 453734
rect 92394 418054 93014 453498
rect 92394 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 93014 418054
rect 92394 417734 93014 417818
rect 92394 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 93014 417734
rect 92394 382054 93014 417498
rect 92394 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 93014 382054
rect 92394 381734 93014 381818
rect 92394 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 93014 381734
rect 92394 346054 93014 381498
rect 92394 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 93014 346054
rect 92394 345734 93014 345818
rect 92394 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 93014 345734
rect 92394 310054 93014 345498
rect 92394 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 93014 310054
rect 92394 309734 93014 309818
rect 92394 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 93014 309734
rect 92394 274054 93014 309498
rect 92394 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 93014 274054
rect 92394 273734 93014 273818
rect 92394 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 93014 273734
rect 92394 238054 93014 273498
rect 92394 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 93014 238054
rect 92394 237734 93014 237818
rect 92394 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 93014 237734
rect 92394 202054 93014 237498
rect 92394 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 93014 202054
rect 92394 201734 93014 201818
rect 92394 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 93014 201734
rect 92394 195244 93014 201498
rect 96114 493774 96734 498064
rect 98502 496909 98562 499530
rect 100894 499530 100988 499590
rect 99834 497494 100454 498064
rect 99834 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 100454 497494
rect 99834 497174 100454 497258
rect 99834 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 100454 497174
rect 98499 496908 98565 496909
rect 98499 496844 98500 496908
rect 98564 496844 98565 496908
rect 98499 496843 98565 496844
rect 96114 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 96734 493774
rect 96114 493454 96734 493538
rect 96114 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 96734 493454
rect 96114 457774 96734 493218
rect 96114 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 96734 457774
rect 96114 457454 96734 457538
rect 96114 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 96734 457454
rect 96114 421774 96734 457218
rect 96114 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 96734 421774
rect 96114 421454 96734 421538
rect 96114 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 96734 421454
rect 96114 385774 96734 421218
rect 96114 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 96734 385774
rect 96114 385454 96734 385538
rect 96114 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 96734 385454
rect 96114 349774 96734 385218
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 96114 313774 96734 349218
rect 96114 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 96734 313774
rect 96114 313454 96734 313538
rect 96114 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 96734 313454
rect 96114 277774 96734 313218
rect 96114 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 96734 277774
rect 96114 277454 96734 277538
rect 96114 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 96734 277454
rect 96114 241774 96734 277218
rect 96114 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 96734 241774
rect 96114 241454 96734 241538
rect 96114 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 96734 241454
rect 96114 205774 96734 241218
rect 96114 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 96734 205774
rect 96114 205454 96734 205538
rect 96114 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 96734 205454
rect 96114 195244 96734 205218
rect 99834 461494 100454 496938
rect 100894 496909 100954 499530
rect 103512 499490 103572 500106
rect 105960 499590 106020 500106
rect 108544 499590 108604 500106
rect 110992 499590 111052 500106
rect 113440 499590 113500 500106
rect 115888 499590 115948 500106
rect 105960 499530 106106 499590
rect 108544 499530 108682 499590
rect 110992 499530 111074 499590
rect 103286 499430 103572 499490
rect 100891 496908 100957 496909
rect 100891 496844 100892 496908
rect 100956 496844 100957 496908
rect 103286 496906 103346 499430
rect 106046 497181 106106 499530
rect 106043 497180 106109 497181
rect 106043 497116 106044 497180
rect 106108 497116 106109 497180
rect 106043 497115 106109 497116
rect 108622 496909 108682 499530
rect 103467 496908 103533 496909
rect 103467 496906 103468 496908
rect 103286 496846 103468 496906
rect 100891 496843 100957 496844
rect 103467 496844 103468 496846
rect 103532 496844 103533 496908
rect 103467 496843 103533 496844
rect 108619 496908 108685 496909
rect 108619 496844 108620 496908
rect 108684 496844 108685 496908
rect 108619 496843 108685 496844
rect 99834 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 100454 461494
rect 99834 461174 100454 461258
rect 99834 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 100454 461174
rect 99834 425494 100454 460938
rect 99834 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 100454 425494
rect 99834 425174 100454 425258
rect 99834 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 100454 425174
rect 99834 389494 100454 424938
rect 99834 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 100454 389494
rect 99834 389174 100454 389258
rect 99834 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 100454 389174
rect 99834 353494 100454 388938
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 99834 317494 100454 352938
rect 99834 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 100454 317494
rect 99834 317174 100454 317258
rect 99834 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 100454 317174
rect 99834 281494 100454 316938
rect 99834 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 100454 281494
rect 99834 281174 100454 281258
rect 99834 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 100454 281174
rect 99834 245494 100454 280938
rect 99834 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 100454 245494
rect 99834 245174 100454 245258
rect 99834 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 100454 245174
rect 99834 209494 100454 244938
rect 99834 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 100454 209494
rect 99834 209174 100454 209258
rect 99834 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 100454 209174
rect 99834 195244 100454 208938
rect 109794 471454 110414 498064
rect 111014 496909 111074 499530
rect 113406 499530 113500 499590
rect 115798 499530 115948 499590
rect 118472 499590 118532 500106
rect 120920 499590 120980 500106
rect 123368 499590 123428 500106
rect 125952 499590 126012 500106
rect 118472 499530 118618 499590
rect 120920 499530 121010 499590
rect 113406 498133 113466 499530
rect 113403 498132 113469 498133
rect 113403 498068 113404 498132
rect 113468 498068 113469 498132
rect 113403 498067 113469 498068
rect 111011 496908 111077 496909
rect 111011 496844 111012 496908
rect 111076 496844 111077 496908
rect 111011 496843 111077 496844
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 195244 110414 218898
rect 113514 475174 114134 497940
rect 115798 496909 115858 499530
rect 115795 496908 115861 496909
rect 115795 496844 115796 496908
rect 115860 496844 115861 496908
rect 115795 496843 115861 496844
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 195244 114134 222618
rect 117234 478894 117854 498064
rect 118558 496909 118618 499530
rect 120950 498133 121010 499530
rect 123342 499530 123428 499590
rect 125918 499530 126012 499590
rect 120947 498132 121013 498133
rect 120947 498068 120948 498132
rect 121012 498068 121013 498132
rect 120947 498067 121013 498068
rect 118555 496908 118621 496909
rect 118555 496844 118556 496908
rect 118620 496844 118621 496908
rect 118555 496843 118621 496844
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 195244 117854 226338
rect 120954 482614 121574 497940
rect 123342 496909 123402 499530
rect 123339 496908 123405 496909
rect 123339 496844 123340 496908
rect 123404 496844 123405 496908
rect 123339 496843 123405 496844
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 195244 121574 230058
rect 124674 486334 125294 498064
rect 125918 496909 125978 499530
rect 125915 496908 125981 496909
rect 125915 496844 125916 496908
rect 125980 496844 125981 496908
rect 125915 496843 125981 496844
rect 124674 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 125294 486334
rect 124674 486014 125294 486098
rect 124674 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 125294 486014
rect 124674 450334 125294 485778
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 124674 414334 125294 449778
rect 124674 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 125294 414334
rect 124674 414014 125294 414098
rect 124674 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 125294 414014
rect 124674 378334 125294 413778
rect 124674 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 125294 378334
rect 124674 378014 125294 378098
rect 124674 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 125294 378014
rect 124674 342334 125294 377778
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 124674 306334 125294 341778
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 124674 270334 125294 305778
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 124674 234334 125294 269778
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 124674 198334 125294 233778
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 124674 195244 125294 197778
rect 128394 490054 129014 498064
rect 128394 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 129014 490054
rect 128394 489734 129014 489818
rect 128394 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 129014 489734
rect 128394 454054 129014 489498
rect 128394 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 129014 454054
rect 128394 453734 129014 453818
rect 128394 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 129014 453734
rect 128394 418054 129014 453498
rect 128394 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 129014 418054
rect 128394 417734 129014 417818
rect 128394 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 129014 417734
rect 128394 382054 129014 417498
rect 128394 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 129014 382054
rect 128394 381734 129014 381818
rect 128394 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 129014 381734
rect 128394 346054 129014 381498
rect 128394 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 129014 346054
rect 128394 345734 129014 345818
rect 128394 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 129014 345734
rect 128394 310054 129014 345498
rect 128394 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 129014 310054
rect 128394 309734 129014 309818
rect 128394 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 129014 309734
rect 128394 274054 129014 309498
rect 128394 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 129014 274054
rect 128394 273734 129014 273818
rect 128394 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 129014 273734
rect 128394 238054 129014 273498
rect 128394 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 129014 238054
rect 128394 237734 129014 237818
rect 128394 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 129014 237734
rect 128394 202054 129014 237498
rect 128394 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 129014 202054
rect 128394 201734 129014 201818
rect 128394 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 129014 201734
rect 128394 195244 129014 201498
rect 132114 493774 132734 498064
rect 132114 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 132734 493774
rect 132114 493454 132734 493538
rect 132114 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 132734 493454
rect 132114 457774 132734 493218
rect 132114 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 132734 457774
rect 132114 457454 132734 457538
rect 132114 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 132734 457454
rect 132114 421774 132734 457218
rect 132114 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 132734 421774
rect 132114 421454 132734 421538
rect 132114 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 132734 421454
rect 132114 385774 132734 421218
rect 132114 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 132734 385774
rect 132114 385454 132734 385538
rect 132114 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 132734 385454
rect 132114 349774 132734 385218
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 132114 313774 132734 349218
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 132114 277774 132734 313218
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 132114 241774 132734 277218
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 132114 205774 132734 241218
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 132114 195244 132734 205218
rect 135834 497494 136454 498064
rect 135834 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 136454 497494
rect 135834 497174 136454 497258
rect 135834 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 136454 497174
rect 135834 461494 136454 496938
rect 135834 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 136454 461494
rect 135834 461174 136454 461258
rect 135834 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 136454 461174
rect 135834 425494 136454 460938
rect 135834 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 136454 425494
rect 135834 425174 136454 425258
rect 135834 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 136454 425174
rect 135834 389494 136454 424938
rect 135834 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 136454 389494
rect 135834 389174 136454 389258
rect 135834 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 136454 389174
rect 135834 353494 136454 388938
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 135834 317494 136454 352938
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 135834 281494 136454 316938
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 135834 245494 136454 280938
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 135834 209494 136454 244938
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 135834 195244 136454 208938
rect 145794 471454 146414 498064
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 195244 146414 218898
rect 149514 475174 150134 498064
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 195244 150134 222618
rect 153234 478894 153854 498064
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 150939 196076 151005 196077
rect 150939 196012 150940 196076
rect 151004 196012 151005 196076
rect 150939 196011 151005 196012
rect 150942 193490 151002 196011
rect 153234 195244 153854 226338
rect 156954 482614 157574 498064
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 195244 157574 230058
rect 160674 486334 161294 521778
rect 160674 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 161294 486334
rect 160674 486014 161294 486098
rect 160674 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 161294 486014
rect 160674 450334 161294 485778
rect 160674 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 161294 450334
rect 160674 450014 161294 450098
rect 160674 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 161294 450014
rect 160674 414334 161294 449778
rect 160674 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 161294 414334
rect 160674 414014 161294 414098
rect 160674 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 161294 414014
rect 160674 378334 161294 413778
rect 160674 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 161294 378334
rect 160674 378014 161294 378098
rect 160674 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 161294 378014
rect 160674 342334 161294 377778
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 160674 306334 161294 341778
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 160674 270334 161294 305778
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 160674 234334 161294 269778
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 150840 193430 151002 193490
rect 150840 193202 150900 193430
rect 20272 187174 20620 187206
rect 20272 186938 20328 187174
rect 20564 186938 20620 187174
rect 20272 186854 20620 186938
rect 20272 186618 20328 186854
rect 20564 186618 20620 186854
rect 20272 186586 20620 186618
rect 156000 187174 156348 187206
rect 156000 186938 156056 187174
rect 156292 186938 156348 187174
rect 156000 186854 156348 186938
rect 156000 186618 156056 186854
rect 156292 186618 156348 186854
rect 156000 186586 156348 186618
rect 20952 183454 21300 183486
rect 20952 183218 21008 183454
rect 21244 183218 21300 183454
rect 20952 183134 21300 183218
rect 20952 182898 21008 183134
rect 21244 182898 21300 183134
rect 20952 182866 21300 182898
rect 155320 183454 155668 183486
rect 155320 183218 155376 183454
rect 155612 183218 155668 183454
rect 155320 183134 155668 183218
rect 155320 182898 155376 183134
rect 155612 182898 155668 183134
rect 155320 182866 155668 182898
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 20272 151174 20620 151206
rect 20272 150938 20328 151174
rect 20564 150938 20620 151174
rect 20272 150854 20620 150938
rect 20272 150618 20328 150854
rect 20564 150618 20620 150854
rect 20272 150586 20620 150618
rect 156000 151174 156348 151206
rect 156000 150938 156056 151174
rect 156292 150938 156348 151174
rect 156000 150854 156348 150938
rect 156000 150618 156056 150854
rect 156292 150618 156348 150854
rect 156000 150586 156348 150618
rect 20952 147454 21300 147486
rect 20952 147218 21008 147454
rect 21244 147218 21300 147454
rect 20952 147134 21300 147218
rect 20952 146898 21008 147134
rect 21244 146898 21300 147134
rect 20952 146866 21300 146898
rect 155320 147454 155668 147486
rect 155320 147218 155376 147454
rect 155612 147218 155668 147454
rect 155320 147134 155668 147218
rect 155320 146898 155376 147134
rect 155612 146898 155668 147134
rect 155320 146866 155668 146898
rect 160674 126334 161294 161778
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 20272 115174 20620 115206
rect 20272 114938 20328 115174
rect 20564 114938 20620 115174
rect 20272 114854 20620 114938
rect 20272 114618 20328 114854
rect 20564 114618 20620 114854
rect 20272 114586 20620 114618
rect 156000 115174 156348 115206
rect 156000 114938 156056 115174
rect 156292 114938 156348 115174
rect 156000 114854 156348 114938
rect 156000 114618 156056 114854
rect 156292 114618 156348 114854
rect 156000 114586 156348 114618
rect 20952 111337 21300 111486
rect 20952 111101 21008 111337
rect 21244 111101 21300 111337
rect 20952 110952 21300 111101
rect 155320 111337 155668 111486
rect 155320 111101 155376 111337
rect 155612 111101 155668 111337
rect 155320 110952 155668 111101
rect 36056 109850 36116 110106
rect 37144 109850 37204 110106
rect 38232 109850 38292 110106
rect 35942 109790 36116 109850
rect 37046 109790 37204 109850
rect 38150 109790 38292 109850
rect 39592 109850 39652 110106
rect 40544 109850 40604 110106
rect 39592 109790 39682 109850
rect 35942 107541 36002 109790
rect 37046 107541 37106 109790
rect 38150 107541 38210 109790
rect 39622 107541 39682 109790
rect 40542 109790 40604 109850
rect 41768 109850 41828 110106
rect 43128 109850 43188 110106
rect 41768 109790 41890 109850
rect 40542 107541 40602 109790
rect 19931 107540 19997 107541
rect 19931 107476 19932 107540
rect 19996 107476 19997 107540
rect 19931 107475 19997 107476
rect 35939 107540 36005 107541
rect 35939 107476 35940 107540
rect 36004 107476 36005 107540
rect 35939 107475 36005 107476
rect 37043 107540 37109 107541
rect 37043 107476 37044 107540
rect 37108 107476 37109 107540
rect 37043 107475 37109 107476
rect 38147 107540 38213 107541
rect 38147 107476 38148 107540
rect 38212 107476 38213 107540
rect 38147 107475 38213 107476
rect 39619 107540 39685 107541
rect 39619 107476 39620 107540
rect 39684 107476 39685 107540
rect 39619 107475 39685 107476
rect 40539 107540 40605 107541
rect 40539 107476 40540 107540
rect 40604 107476 40605 107540
rect 40539 107475 40605 107476
rect 41830 107405 41890 109790
rect 43118 109790 43188 109850
rect 44216 109850 44276 110106
rect 45440 109850 45500 110106
rect 44216 109790 44282 109850
rect 43118 107541 43178 109790
rect 44222 107541 44282 109790
rect 45326 109790 45500 109850
rect 46528 109850 46588 110106
rect 47616 109850 47676 110106
rect 48296 109850 48356 110106
rect 48704 109850 48764 110106
rect 46528 109790 46674 109850
rect 45326 107541 45386 109790
rect 46614 107541 46674 109790
rect 47534 109790 47676 109850
rect 48270 109790 48356 109850
rect 48638 109790 48764 109850
rect 50064 109850 50124 110106
rect 50064 109790 50170 109850
rect 47534 107541 47594 109790
rect 48270 109037 48330 109790
rect 48267 109036 48333 109037
rect 48267 108972 48268 109036
rect 48332 108972 48333 109036
rect 48267 108971 48333 108972
rect 48638 107541 48698 109790
rect 50110 107541 50170 109790
rect 50744 109581 50804 110106
rect 51288 109850 51348 110106
rect 52376 109850 52436 110106
rect 53464 109850 53524 110106
rect 51214 109790 51348 109850
rect 52318 109790 52436 109850
rect 53422 109790 53524 109850
rect 53600 109850 53660 110106
rect 54552 109850 54612 110106
rect 55912 109850 55972 110106
rect 53600 109790 53666 109850
rect 50741 109580 50807 109581
rect 50741 109516 50742 109580
rect 50806 109516 50807 109580
rect 50741 109515 50807 109516
rect 51214 107541 51274 109790
rect 52318 107541 52378 109790
rect 53422 107541 53482 109790
rect 53606 108765 53666 109790
rect 54526 109790 54612 109850
rect 55814 109790 55972 109850
rect 53603 108764 53669 108765
rect 53603 108700 53604 108764
rect 53668 108700 53669 108764
rect 53603 108699 53669 108700
rect 43115 107540 43181 107541
rect 43115 107476 43116 107540
rect 43180 107476 43181 107540
rect 43115 107475 43181 107476
rect 44219 107540 44285 107541
rect 44219 107476 44220 107540
rect 44284 107476 44285 107540
rect 44219 107475 44285 107476
rect 45323 107540 45389 107541
rect 45323 107476 45324 107540
rect 45388 107476 45389 107540
rect 45323 107475 45389 107476
rect 46611 107540 46677 107541
rect 46611 107476 46612 107540
rect 46676 107476 46677 107540
rect 46611 107475 46677 107476
rect 47531 107540 47597 107541
rect 47531 107476 47532 107540
rect 47596 107476 47597 107540
rect 47531 107475 47597 107476
rect 48635 107540 48701 107541
rect 48635 107476 48636 107540
rect 48700 107476 48701 107540
rect 48635 107475 48701 107476
rect 50107 107540 50173 107541
rect 50107 107476 50108 107540
rect 50172 107476 50173 107540
rect 50107 107475 50173 107476
rect 51211 107540 51277 107541
rect 51211 107476 51212 107540
rect 51276 107476 51277 107540
rect 51211 107475 51277 107476
rect 52315 107540 52381 107541
rect 52315 107476 52316 107540
rect 52380 107476 52381 107540
rect 52315 107475 52381 107476
rect 53419 107540 53485 107541
rect 53419 107476 53420 107540
rect 53484 107476 53485 107540
rect 53419 107475 53485 107476
rect 41827 107404 41893 107405
rect 41827 107340 41828 107404
rect 41892 107340 41893 107404
rect 41827 107339 41893 107340
rect 54526 107133 54586 109790
rect 55814 107133 55874 109790
rect 56048 109581 56108 110106
rect 57000 109850 57060 110106
rect 58088 109850 58148 110106
rect 57000 109790 57162 109850
rect 56045 109580 56111 109581
rect 56045 109516 56046 109580
rect 56110 109516 56111 109580
rect 56045 109515 56111 109516
rect 57102 107405 57162 109790
rect 58022 109790 58148 109850
rect 58496 109850 58556 110106
rect 59448 109850 59508 110106
rect 60672 109850 60732 110106
rect 58496 109790 58634 109850
rect 59448 109790 59554 109850
rect 57099 107404 57165 107405
rect 57099 107340 57100 107404
rect 57164 107340 57165 107404
rect 57099 107339 57165 107340
rect 54523 107132 54589 107133
rect 54523 107068 54524 107132
rect 54588 107068 54589 107132
rect 54523 107067 54589 107068
rect 55811 107132 55877 107133
rect 55811 107068 55812 107132
rect 55876 107068 55877 107132
rect 55811 107067 55877 107068
rect 57102 106317 57162 107339
rect 58022 107269 58082 109790
rect 58019 107268 58085 107269
rect 58019 107204 58020 107268
rect 58084 107204 58085 107268
rect 58019 107203 58085 107204
rect 58574 106725 58634 109790
rect 59494 107541 59554 109790
rect 60598 109790 60732 109850
rect 60598 107541 60658 109790
rect 61080 109581 61140 110106
rect 61760 109850 61820 110106
rect 62848 109850 62908 110106
rect 61702 109790 61820 109850
rect 62806 109790 62908 109850
rect 63528 109850 63588 110106
rect 63936 109850 63996 110106
rect 65296 109850 65356 110106
rect 65976 109850 66036 110106
rect 66384 109850 66444 110106
rect 67608 109850 67668 110106
rect 63528 109790 63602 109850
rect 61077 109580 61143 109581
rect 61077 109516 61078 109580
rect 61142 109516 61143 109580
rect 61077 109515 61143 109516
rect 61702 107541 61762 109790
rect 62806 107541 62866 109790
rect 63542 107541 63602 109790
rect 63910 109790 63996 109850
rect 65198 109790 65356 109850
rect 65934 109790 66036 109850
rect 66302 109790 66444 109850
rect 67590 109790 67668 109850
rect 68288 109850 68348 110106
rect 68696 109850 68756 110106
rect 68288 109790 68386 109850
rect 63910 107541 63970 109790
rect 65198 107541 65258 109790
rect 65934 108901 65994 109790
rect 65931 108900 65997 108901
rect 65931 108836 65932 108900
rect 65996 108836 65997 108900
rect 65931 108835 65997 108836
rect 66302 107541 66362 109790
rect 67590 107541 67650 109790
rect 68326 109037 68386 109790
rect 68694 109790 68756 109850
rect 69784 109850 69844 110106
rect 71008 109850 71068 110106
rect 69784 109790 69858 109850
rect 68323 109036 68389 109037
rect 68323 108972 68324 109036
rect 68388 108972 68389 109036
rect 68323 108971 68389 108972
rect 68694 107541 68754 109790
rect 69798 107541 69858 109790
rect 70902 109790 71068 109850
rect 71144 109850 71204 110106
rect 72232 109850 72292 110106
rect 73320 109850 73380 110106
rect 71144 109790 71330 109850
rect 59491 107540 59557 107541
rect 59491 107476 59492 107540
rect 59556 107476 59557 107540
rect 59491 107475 59557 107476
rect 60595 107540 60661 107541
rect 60595 107476 60596 107540
rect 60660 107476 60661 107540
rect 60595 107475 60661 107476
rect 61699 107540 61765 107541
rect 61699 107476 61700 107540
rect 61764 107476 61765 107540
rect 61699 107475 61765 107476
rect 62803 107540 62869 107541
rect 62803 107476 62804 107540
rect 62868 107476 62869 107540
rect 62803 107475 62869 107476
rect 63539 107540 63605 107541
rect 63539 107476 63540 107540
rect 63604 107476 63605 107540
rect 63539 107475 63605 107476
rect 63907 107540 63973 107541
rect 63907 107476 63908 107540
rect 63972 107476 63973 107540
rect 63907 107475 63973 107476
rect 65195 107540 65261 107541
rect 65195 107476 65196 107540
rect 65260 107476 65261 107540
rect 65195 107475 65261 107476
rect 66299 107540 66365 107541
rect 66299 107476 66300 107540
rect 66364 107476 66365 107540
rect 66299 107475 66365 107476
rect 67587 107540 67653 107541
rect 67587 107476 67588 107540
rect 67652 107476 67653 107540
rect 67587 107475 67653 107476
rect 68691 107540 68757 107541
rect 68691 107476 68692 107540
rect 68756 107476 68757 107540
rect 68691 107475 68757 107476
rect 69795 107540 69861 107541
rect 69795 107476 69796 107540
rect 69860 107476 69861 107540
rect 69795 107475 69861 107476
rect 70902 107405 70962 109790
rect 71270 107541 71330 109790
rect 72190 109790 72292 109850
rect 73294 109790 73380 109850
rect 73592 109850 73652 110106
rect 74408 109850 74468 110106
rect 75768 109850 75828 110106
rect 73592 109790 73722 109850
rect 72190 107541 72250 109790
rect 73294 107541 73354 109790
rect 73662 107541 73722 109790
rect 74398 109790 74468 109850
rect 75686 109790 75828 109850
rect 76040 109850 76100 110106
rect 76992 109850 77052 110106
rect 78080 109850 78140 110106
rect 78488 109850 78548 110106
rect 76040 109790 76114 109850
rect 74398 107541 74458 109790
rect 75686 107541 75746 109790
rect 76054 107541 76114 109790
rect 76974 109790 77052 109850
rect 78078 109790 78140 109850
rect 78446 109790 78548 109850
rect 79168 109850 79228 110106
rect 80936 109850 80996 110106
rect 83520 109850 83580 110106
rect 85968 109850 86028 110106
rect 88280 109850 88340 110106
rect 91000 109850 91060 110106
rect 79168 109790 79242 109850
rect 80936 109790 81082 109850
rect 83520 109790 83658 109850
rect 85968 109790 86050 109850
rect 71267 107540 71333 107541
rect 71267 107476 71268 107540
rect 71332 107476 71333 107540
rect 71267 107475 71333 107476
rect 72187 107540 72253 107541
rect 72187 107476 72188 107540
rect 72252 107476 72253 107540
rect 72187 107475 72253 107476
rect 73291 107540 73357 107541
rect 73291 107476 73292 107540
rect 73356 107476 73357 107540
rect 73291 107475 73357 107476
rect 73659 107540 73725 107541
rect 73659 107476 73660 107540
rect 73724 107476 73725 107540
rect 73659 107475 73725 107476
rect 74395 107540 74461 107541
rect 74395 107476 74396 107540
rect 74460 107476 74461 107540
rect 74395 107475 74461 107476
rect 75683 107540 75749 107541
rect 75683 107476 75684 107540
rect 75748 107476 75749 107540
rect 75683 107475 75749 107476
rect 76051 107540 76117 107541
rect 76051 107476 76052 107540
rect 76116 107476 76117 107540
rect 76051 107475 76117 107476
rect 70899 107404 70965 107405
rect 70899 107340 70900 107404
rect 70964 107340 70965 107404
rect 70899 107339 70965 107340
rect 76974 107269 77034 109790
rect 78078 107541 78138 109790
rect 78446 107541 78506 109790
rect 79182 107541 79242 109790
rect 78075 107540 78141 107541
rect 78075 107476 78076 107540
rect 78140 107476 78141 107540
rect 78075 107475 78141 107476
rect 78443 107540 78509 107541
rect 78443 107476 78444 107540
rect 78508 107476 78509 107540
rect 78443 107475 78509 107476
rect 79179 107540 79245 107541
rect 79179 107476 79180 107540
rect 79244 107476 79245 107540
rect 79179 107475 79245 107476
rect 81022 107269 81082 109790
rect 76971 107268 77037 107269
rect 76971 107204 76972 107268
rect 77036 107204 77037 107268
rect 76971 107203 77037 107204
rect 81019 107268 81085 107269
rect 81019 107204 81020 107268
rect 81084 107204 81085 107268
rect 81019 107203 81085 107204
rect 83598 107133 83658 109790
rect 85990 107541 86050 109790
rect 88198 109790 88340 109850
rect 90958 109790 91060 109850
rect 93448 109850 93508 110106
rect 95896 109850 95956 110106
rect 98480 109850 98540 110106
rect 100928 109850 100988 110106
rect 103512 109850 103572 110106
rect 93448 109790 93594 109850
rect 95896 109790 95986 109850
rect 98480 109790 98562 109850
rect 88198 107541 88258 109790
rect 90958 108765 91018 109790
rect 90955 108764 91021 108765
rect 90955 108700 90956 108764
rect 91020 108700 91021 108764
rect 90955 108699 91021 108700
rect 93534 107541 93594 109790
rect 95926 108629 95986 109790
rect 95923 108628 95989 108629
rect 95923 108564 95924 108628
rect 95988 108564 95989 108628
rect 95923 108563 95989 108564
rect 98502 107541 98562 109790
rect 100894 109790 100988 109850
rect 103286 109790 103572 109850
rect 100894 109037 100954 109790
rect 100891 109036 100957 109037
rect 100891 108972 100892 109036
rect 100956 108972 100957 109036
rect 100891 108971 100957 108972
rect 85987 107540 86053 107541
rect 85987 107476 85988 107540
rect 86052 107476 86053 107540
rect 85987 107475 86053 107476
rect 88195 107540 88261 107541
rect 88195 107476 88196 107540
rect 88260 107476 88261 107540
rect 88195 107475 88261 107476
rect 93531 107540 93597 107541
rect 93531 107476 93532 107540
rect 93596 107476 93597 107540
rect 93531 107475 93597 107476
rect 98499 107540 98565 107541
rect 98499 107476 98500 107540
rect 98564 107476 98565 107540
rect 98499 107475 98565 107476
rect 83595 107132 83661 107133
rect 83595 107068 83596 107132
rect 83660 107068 83661 107132
rect 103286 107130 103346 109790
rect 105960 109581 106020 110106
rect 108544 109581 108604 110106
rect 110992 109850 111052 110106
rect 113440 109850 113500 110106
rect 115888 109850 115948 110106
rect 110992 109790 111074 109850
rect 105957 109580 106023 109581
rect 105957 109516 105958 109580
rect 106022 109516 106023 109580
rect 105957 109515 106023 109516
rect 108541 109580 108607 109581
rect 108541 109516 108542 109580
rect 108606 109516 108607 109580
rect 108541 109515 108607 109516
rect 111014 109037 111074 109790
rect 113406 109790 113500 109850
rect 115798 109790 115948 109850
rect 118472 109850 118532 110106
rect 120920 109850 120980 110106
rect 123368 109850 123428 110106
rect 125952 109850 126012 110106
rect 118472 109790 118618 109850
rect 120920 109790 121010 109850
rect 113406 109037 113466 109790
rect 111011 109036 111077 109037
rect 111011 108972 111012 109036
rect 111076 108972 111077 109036
rect 111011 108971 111077 108972
rect 113403 109036 113469 109037
rect 113403 108972 113404 109036
rect 113468 108972 113469 109036
rect 113403 108971 113469 108972
rect 103286 107070 103530 107130
rect 83595 107067 83661 107068
rect 103470 106997 103530 107070
rect 103467 106996 103533 106997
rect 103467 106932 103468 106996
rect 103532 106932 103533 106996
rect 103467 106931 103533 106932
rect 115798 106861 115858 109790
rect 118558 108493 118618 109790
rect 118555 108492 118621 108493
rect 118555 108428 118556 108492
rect 118620 108428 118621 108492
rect 118555 108427 118621 108428
rect 120950 107541 121010 109790
rect 123342 109790 123428 109850
rect 125918 109790 126012 109850
rect 123342 107541 123402 109790
rect 125918 109037 125978 109790
rect 125915 109036 125981 109037
rect 125915 108972 125916 109036
rect 125980 108972 125981 109036
rect 125915 108971 125981 108972
rect 120947 107540 121013 107541
rect 120947 107476 120948 107540
rect 121012 107476 121013 107540
rect 120947 107475 121013 107476
rect 123339 107540 123405 107541
rect 123339 107476 123340 107540
rect 123404 107476 123405 107540
rect 123339 107475 123405 107476
rect 115795 106860 115861 106861
rect 115795 106796 115796 106860
rect 115860 106796 115861 106860
rect 115795 106795 115861 106796
rect 58571 106724 58637 106725
rect 58571 106660 58572 106724
rect 58636 106660 58637 106724
rect 58571 106659 58637 106660
rect 57099 106316 57165 106317
rect 57099 106252 57100 106316
rect 57164 106252 57165 106316
rect 57099 106251 57165 106252
rect 150755 105364 150821 105365
rect 150755 105300 150756 105364
rect 150820 105300 150821 105364
rect 150755 105299 150821 105300
rect 150758 103530 150818 105299
rect 150758 103470 150900 103530
rect 150840 103202 150900 103470
rect 160674 90334 161294 125778
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 20272 79174 20620 79206
rect 20272 78938 20328 79174
rect 20564 78938 20620 79174
rect 20272 78854 20620 78938
rect 20272 78618 20328 78854
rect 20564 78618 20620 78854
rect 20272 78586 20620 78618
rect 156000 79174 156348 79206
rect 156000 78938 156056 79174
rect 156292 78938 156348 79174
rect 156000 78854 156348 78938
rect 156000 78618 156056 78854
rect 156292 78618 156348 78854
rect 156000 78586 156348 78618
rect 20952 75454 21300 75486
rect 20952 75218 21008 75454
rect 21244 75218 21300 75454
rect 20952 75134 21300 75218
rect 20952 74898 21008 75134
rect 21244 74898 21300 75134
rect 20952 74866 21300 74898
rect 155320 75454 155668 75486
rect 155320 75218 155376 75454
rect 155612 75218 155668 75454
rect 155320 75134 155668 75218
rect 155320 74898 155376 75134
rect 155612 74898 155668 75134
rect 155320 74866 155668 74898
rect 160674 54334 161294 89778
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 20272 43174 20620 43206
rect 20272 42938 20328 43174
rect 20564 42938 20620 43174
rect 20272 42854 20620 42938
rect 20272 42618 20328 42854
rect 20564 42618 20620 42854
rect 20272 42586 20620 42618
rect 156000 43174 156348 43206
rect 156000 42938 156056 43174
rect 156292 42938 156348 43174
rect 156000 42854 156348 42938
rect 156000 42618 156056 42854
rect 156292 42618 156348 42854
rect 156000 42586 156348 42618
rect 20952 39454 21300 39486
rect 20952 39218 21008 39454
rect 21244 39218 21300 39454
rect 20952 39134 21300 39218
rect 20952 38898 21008 39134
rect 21244 38898 21300 39134
rect 20952 38866 21300 38898
rect 155320 39454 155668 39486
rect 155320 39218 155376 39454
rect 155612 39218 155668 39454
rect 155320 39134 155668 39218
rect 155320 38898 155376 39134
rect 155612 38898 155668 39134
rect 155320 38866 155668 38898
rect 19195 28116 19261 28117
rect 19195 28052 19196 28116
rect 19260 28052 19261 28116
rect 19195 28051 19261 28052
rect 36056 19410 36116 20060
rect 37144 19410 37204 20060
rect 35942 19350 36116 19410
rect 37046 19350 37204 19410
rect 38232 19410 38292 20060
rect 39592 19410 39652 20060
rect 40544 19410 40604 20060
rect 41768 19410 41828 20060
rect 43128 19410 43188 20060
rect 38232 19350 38578 19410
rect 39592 19350 39682 19410
rect 16674 -4186 17294 17778
rect 19011 17780 19077 17781
rect 19011 17716 19012 17780
rect 19076 17716 19077 17780
rect 19011 17715 19077 17716
rect 35942 17237 36002 19350
rect 37046 17917 37106 19350
rect 37043 17916 37109 17917
rect 37043 17852 37044 17916
rect 37108 17852 37109 17916
rect 37043 17851 37109 17852
rect 35939 17236 36005 17237
rect 35939 17172 35940 17236
rect 36004 17172 36005 17236
rect 35939 17171 36005 17172
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 37794 3454 38414 17940
rect 38518 17509 38578 19350
rect 38515 17508 38581 17509
rect 38515 17444 38516 17508
rect 38580 17444 38581 17508
rect 38515 17443 38581 17444
rect 39622 17237 39682 19350
rect 40542 19350 40604 19410
rect 41646 19350 41828 19410
rect 43118 19350 43188 19410
rect 44216 19410 44276 20060
rect 45440 19410 45500 20060
rect 44216 19350 44282 19410
rect 40542 17645 40602 19350
rect 41646 18189 41706 19350
rect 41643 18188 41709 18189
rect 41643 18124 41644 18188
rect 41708 18124 41709 18188
rect 41643 18123 41709 18124
rect 40539 17644 40605 17645
rect 40539 17580 40540 17644
rect 40604 17580 40605 17644
rect 40539 17579 40605 17580
rect 39619 17236 39685 17237
rect 39619 17172 39620 17236
rect 39684 17172 39685 17236
rect 39619 17171 39685 17172
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 7174 42134 17940
rect 43118 17917 43178 19350
rect 44222 17917 44282 19350
rect 45326 19350 45500 19410
rect 46528 19410 46588 20060
rect 47616 19410 47676 20060
rect 48296 19410 48356 20060
rect 48704 19410 48764 20060
rect 46528 19350 46674 19410
rect 45326 18189 45386 19350
rect 45323 18188 45389 18189
rect 45323 18124 45324 18188
rect 45388 18124 45389 18188
rect 45323 18123 45389 18124
rect 43115 17916 43181 17917
rect 43115 17852 43116 17916
rect 43180 17852 43181 17916
rect 43115 17851 43181 17852
rect 44219 17916 44285 17917
rect 44219 17852 44220 17916
rect 44284 17852 44285 17916
rect 44219 17851 44285 17852
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 10894 45854 17940
rect 46614 17917 46674 19350
rect 47534 19350 47676 19410
rect 48270 19350 48356 19410
rect 48638 19350 48764 19410
rect 50064 19410 50124 20060
rect 50744 19410 50804 20060
rect 51288 19410 51348 20060
rect 52376 19549 52436 20060
rect 53464 19549 53524 20060
rect 52373 19548 52439 19549
rect 52373 19484 52374 19548
rect 52438 19484 52439 19548
rect 52373 19483 52439 19484
rect 53461 19548 53527 19549
rect 53461 19484 53462 19548
rect 53526 19484 53527 19548
rect 53461 19483 53527 19484
rect 53600 19410 53660 20060
rect 54552 19410 54612 20060
rect 55912 19549 55972 20060
rect 55909 19548 55975 19549
rect 55909 19484 55910 19548
rect 55974 19484 55975 19548
rect 55909 19483 55975 19484
rect 56048 19410 56108 20060
rect 57000 19410 57060 20060
rect 50064 19350 50170 19410
rect 50744 19350 50906 19410
rect 51288 19350 51458 19410
rect 53600 19350 53666 19410
rect 47534 17917 47594 19350
rect 46611 17916 46677 17917
rect 46611 17852 46612 17916
rect 46676 17852 46677 17916
rect 46611 17851 46677 17852
rect 47531 17916 47597 17917
rect 47531 17852 47532 17916
rect 47596 17852 47597 17916
rect 47531 17851 47597 17852
rect 48270 17781 48330 19350
rect 48638 17917 48698 19350
rect 48635 17916 48701 17917
rect 48635 17852 48636 17916
rect 48700 17852 48701 17916
rect 48635 17851 48701 17852
rect 48267 17780 48333 17781
rect 48267 17716 48268 17780
rect 48332 17716 48333 17780
rect 48267 17715 48333 17716
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 18064
rect 50110 17917 50170 19350
rect 50846 18733 50906 19350
rect 50843 18732 50909 18733
rect 50843 18668 50844 18732
rect 50908 18668 50909 18732
rect 50843 18667 50909 18668
rect 51398 17917 51458 19350
rect 53606 18733 53666 19350
rect 54526 19350 54612 19410
rect 55998 19350 56108 19410
rect 56918 19350 57060 19410
rect 58088 19410 58148 20060
rect 58496 19410 58556 20060
rect 59448 19410 59508 20060
rect 60672 19410 60732 20060
rect 58088 19350 58266 19410
rect 58496 19350 58634 19410
rect 59448 19350 59554 19410
rect 53603 18732 53669 18733
rect 53603 18668 53604 18732
rect 53668 18668 53669 18732
rect 53603 18667 53669 18668
rect 52674 18023 53294 18064
rect 50107 17916 50173 17917
rect 50107 17852 50108 17916
rect 50172 17852 50173 17916
rect 50107 17851 50173 17852
rect 51395 17916 51461 17917
rect 51395 17852 51396 17916
rect 51460 17852 51461 17916
rect 51395 17851 51461 17852
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 17787 52706 18023
rect 52942 17787 53026 18023
rect 53262 17787 53294 18023
rect 52674 -4186 53294 17787
rect 54526 17645 54586 19350
rect 55998 18869 56058 19350
rect 55995 18868 56061 18869
rect 55995 18804 55996 18868
rect 56060 18804 56061 18868
rect 55995 18803 56061 18804
rect 54523 17644 54589 17645
rect 54523 17580 54524 17644
rect 54588 17580 54589 17644
rect 54523 17579 54589 17580
rect 56918 17373 56978 19350
rect 58206 18869 58266 19350
rect 58203 18868 58269 18869
rect 58203 18804 58204 18868
rect 58268 18804 58269 18868
rect 58203 18803 58269 18804
rect 58206 17509 58266 18803
rect 58203 17508 58269 17509
rect 58203 17444 58204 17508
rect 58268 17444 58269 17508
rect 58203 17443 58269 17444
rect 56915 17372 56981 17373
rect 56915 17308 56916 17372
rect 56980 17308 56981 17372
rect 56915 17307 56981 17308
rect 58574 17101 58634 19350
rect 59494 17917 59554 19350
rect 60598 19350 60732 19410
rect 61080 19410 61140 20060
rect 61760 19410 61820 20060
rect 62848 19410 62908 20060
rect 61080 19350 61210 19410
rect 60598 17917 60658 19350
rect 61150 17917 61210 19350
rect 61702 19350 61820 19410
rect 62806 19350 62908 19410
rect 63528 19410 63588 20060
rect 63936 19410 63996 20060
rect 65296 19410 65356 20060
rect 65976 19410 66036 20060
rect 66384 19410 66444 20060
rect 67608 19410 67668 20060
rect 63528 19350 63602 19410
rect 59491 17916 59557 17917
rect 59491 17852 59492 17916
rect 59556 17852 59557 17916
rect 59491 17851 59557 17852
rect 60595 17916 60661 17917
rect 60595 17852 60596 17916
rect 60660 17852 60661 17916
rect 60595 17851 60661 17852
rect 61147 17916 61213 17917
rect 61147 17852 61148 17916
rect 61212 17852 61213 17916
rect 61147 17851 61213 17852
rect 61702 17237 61762 19350
rect 62806 17237 62866 19350
rect 63542 17917 63602 19350
rect 63910 19350 63996 19410
rect 65198 19350 65356 19410
rect 65934 19350 66036 19410
rect 66302 19350 66444 19410
rect 67590 19350 67668 19410
rect 68288 19410 68348 20060
rect 68696 19410 68756 20060
rect 68288 19350 68386 19410
rect 63539 17916 63605 17917
rect 63539 17852 63540 17916
rect 63604 17852 63605 17916
rect 63539 17851 63605 17852
rect 63910 17237 63970 19350
rect 65198 17373 65258 19350
rect 65934 17917 65994 19350
rect 65931 17916 65997 17917
rect 65931 17852 65932 17916
rect 65996 17852 65997 17916
rect 65931 17851 65997 17852
rect 66302 17373 66362 19350
rect 67590 17373 67650 19350
rect 68326 17645 68386 19350
rect 68694 19350 68756 19410
rect 69784 19410 69844 20060
rect 71008 19410 71068 20060
rect 69784 19350 69858 19410
rect 68694 17917 68754 19350
rect 68691 17916 68757 17917
rect 68691 17852 68692 17916
rect 68756 17852 68757 17916
rect 68691 17851 68757 17852
rect 68323 17644 68389 17645
rect 68323 17580 68324 17644
rect 68388 17580 68389 17644
rect 68323 17579 68389 17580
rect 65195 17372 65261 17373
rect 65195 17308 65196 17372
rect 65260 17308 65261 17372
rect 65195 17307 65261 17308
rect 66299 17372 66365 17373
rect 66299 17308 66300 17372
rect 66364 17308 66365 17372
rect 66299 17307 66365 17308
rect 67587 17372 67653 17373
rect 67587 17308 67588 17372
rect 67652 17308 67653 17372
rect 67587 17307 67653 17308
rect 69798 17237 69858 19350
rect 70902 19350 71068 19410
rect 71144 19410 71204 20060
rect 72232 19410 72292 20060
rect 73320 19410 73380 20060
rect 71144 19350 71330 19410
rect 70902 17237 70962 19350
rect 71270 17645 71330 19350
rect 72190 19350 72292 19410
rect 73294 19350 73380 19410
rect 73592 19410 73652 20060
rect 74408 19410 74468 20060
rect 75768 19410 75828 20060
rect 73592 19350 73722 19410
rect 72190 17917 72250 19350
rect 72187 17916 72253 17917
rect 72187 17852 72188 17916
rect 72252 17852 72253 17916
rect 72187 17851 72253 17852
rect 71267 17644 71333 17645
rect 71267 17580 71268 17644
rect 71332 17580 71333 17644
rect 71267 17579 71333 17580
rect 73294 17373 73354 19350
rect 73662 18869 73722 19350
rect 74398 19350 74468 19410
rect 75686 19350 75828 19410
rect 76040 19410 76100 20060
rect 76992 19410 77052 20060
rect 76040 19350 76114 19410
rect 73659 18868 73725 18869
rect 73659 18804 73660 18868
rect 73724 18804 73725 18868
rect 73659 18803 73725 18804
rect 74398 18189 74458 19350
rect 74395 18188 74461 18189
rect 74395 18124 74396 18188
rect 74460 18124 74461 18188
rect 74395 18123 74461 18124
rect 73291 17372 73357 17373
rect 73291 17308 73292 17372
rect 73356 17308 73357 17372
rect 73291 17307 73357 17308
rect 61699 17236 61765 17237
rect 61699 17172 61700 17236
rect 61764 17172 61765 17236
rect 61699 17171 61765 17172
rect 62803 17236 62869 17237
rect 62803 17172 62804 17236
rect 62868 17172 62869 17236
rect 62803 17171 62869 17172
rect 63907 17236 63973 17237
rect 63907 17172 63908 17236
rect 63972 17172 63973 17236
rect 63907 17171 63973 17172
rect 69795 17236 69861 17237
rect 69795 17172 69796 17236
rect 69860 17172 69861 17236
rect 69795 17171 69861 17172
rect 70899 17236 70965 17237
rect 70899 17172 70900 17236
rect 70964 17172 70965 17236
rect 70899 17171 70965 17172
rect 58571 17100 58637 17101
rect 58571 17036 58572 17100
rect 58636 17036 58637 17100
rect 58571 17035 58637 17036
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 73794 3454 74414 17940
rect 75686 17237 75746 19350
rect 76054 19005 76114 19350
rect 76974 19350 77052 19410
rect 78080 19410 78140 20060
rect 78488 19410 78548 20060
rect 78080 19350 78322 19410
rect 76051 19004 76117 19005
rect 76051 18940 76052 19004
rect 76116 18940 76117 19004
rect 76051 18939 76117 18940
rect 76974 17509 77034 19350
rect 76971 17508 77037 17509
rect 76971 17444 76972 17508
rect 77036 17444 77037 17508
rect 76971 17443 77037 17444
rect 75683 17236 75749 17237
rect 75683 17172 75684 17236
rect 75748 17172 75749 17236
rect 75683 17171 75749 17172
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 7174 78134 17940
rect 78262 16965 78322 19350
rect 78446 19350 78548 19410
rect 79168 19410 79228 20060
rect 80936 19410 80996 20060
rect 83520 19410 83580 20060
rect 85968 19410 86028 20060
rect 88280 19410 88340 20060
rect 91000 19410 91060 20060
rect 79168 19350 79242 19410
rect 80936 19350 81082 19410
rect 83520 19350 83658 19410
rect 85968 19350 86050 19410
rect 78446 17917 78506 19350
rect 78443 17916 78509 17917
rect 78443 17852 78444 17916
rect 78508 17852 78509 17916
rect 78443 17851 78509 17852
rect 79182 17509 79242 19350
rect 81022 19005 81082 19350
rect 81019 19004 81085 19005
rect 81019 18940 81020 19004
rect 81084 18940 81085 19004
rect 81019 18939 81085 18940
rect 79179 17508 79245 17509
rect 79179 17444 79180 17508
rect 79244 17444 79245 17508
rect 79179 17443 79245 17444
rect 78259 16964 78325 16965
rect 78259 16900 78260 16964
rect 78324 16900 78325 16964
rect 78259 16899 78325 16900
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 10894 81854 18064
rect 83598 17645 83658 19350
rect 85990 19141 86050 19350
rect 88198 19350 88340 19410
rect 90958 19350 91060 19410
rect 93448 19410 93508 20060
rect 95896 19410 95956 20060
rect 98480 19410 98540 20060
rect 100928 19410 100988 20060
rect 93448 19350 93594 19410
rect 95896 19350 95986 19410
rect 98480 19350 98562 19410
rect 85987 19140 86053 19141
rect 85987 19076 85988 19140
rect 86052 19076 86053 19140
rect 85987 19075 86053 19076
rect 83595 17644 83661 17645
rect 83595 17580 83596 17644
rect 83660 17580 83661 17644
rect 83595 17579 83661 17580
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 18064
rect 88198 17509 88258 19350
rect 90958 19141 91018 19350
rect 90955 19140 91021 19141
rect 90955 19076 90956 19140
rect 91020 19076 91021 19140
rect 90955 19075 91021 19076
rect 88674 18023 89294 18064
rect 88674 17787 88706 18023
rect 88942 17787 89026 18023
rect 89262 17787 89294 18023
rect 88195 17508 88261 17509
rect 88195 17444 88196 17508
rect 88260 17444 88261 17508
rect 88195 17443 88261 17444
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 -4186 89294 17787
rect 93534 17509 93594 19350
rect 95926 19277 95986 19350
rect 95923 19276 95989 19277
rect 95923 19212 95924 19276
rect 95988 19212 95989 19276
rect 95923 19211 95989 19212
rect 93531 17508 93597 17509
rect 93531 17444 93532 17508
rect 93596 17444 93597 17508
rect 93531 17443 93597 17444
rect 98502 17373 98562 19350
rect 100894 19350 100988 19410
rect 103512 19410 103572 20060
rect 105960 19410 106020 20060
rect 108544 19410 108604 20060
rect 110992 19410 111052 20060
rect 113440 19410 113500 20060
rect 115888 19410 115948 20060
rect 103512 19350 103714 19410
rect 105960 19350 106106 19410
rect 108544 19350 108682 19410
rect 110992 19350 111074 19410
rect 100894 19277 100954 19350
rect 103654 19277 103714 19350
rect 100891 19276 100957 19277
rect 100891 19212 100892 19276
rect 100956 19212 100957 19276
rect 100891 19211 100957 19212
rect 103651 19276 103717 19277
rect 103651 19212 103652 19276
rect 103716 19212 103717 19276
rect 103651 19211 103717 19212
rect 106046 18597 106106 19350
rect 108622 18597 108682 19350
rect 106043 18596 106109 18597
rect 106043 18532 106044 18596
rect 106108 18532 106109 18596
rect 106043 18531 106109 18532
rect 108619 18596 108685 18597
rect 108619 18532 108620 18596
rect 108684 18532 108685 18596
rect 108619 18531 108685 18532
rect 98499 17372 98565 17373
rect 98499 17308 98500 17372
rect 98564 17308 98565 17372
rect 98499 17307 98565 17308
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 109794 3454 110414 18064
rect 111014 17373 111074 19350
rect 113406 19350 113500 19410
rect 115798 19350 115948 19410
rect 118472 19410 118532 20060
rect 120920 19410 120980 20060
rect 123368 19410 123428 20060
rect 125952 19410 126012 20060
rect 118472 19350 118618 19410
rect 120920 19350 121010 19410
rect 113406 18461 113466 19350
rect 113403 18460 113469 18461
rect 113403 18396 113404 18460
rect 113468 18396 113469 18460
rect 113403 18395 113469 18396
rect 111011 17372 111077 17373
rect 111011 17308 111012 17372
rect 111076 17308 111077 17372
rect 111011 17307 111077 17308
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 7174 114134 17940
rect 115798 17645 115858 19350
rect 118558 19277 118618 19350
rect 118555 19276 118621 19277
rect 118555 19212 118556 19276
rect 118620 19212 118621 19276
rect 118555 19211 118621 19212
rect 120950 19141 121010 19350
rect 122606 19350 123428 19410
rect 125918 19350 126012 19410
rect 120947 19140 121013 19141
rect 120947 19076 120948 19140
rect 121012 19076 121013 19140
rect 120947 19075 121013 19076
rect 115795 17644 115861 17645
rect 115795 17580 115796 17644
rect 115860 17580 115861 17644
rect 115795 17579 115861 17580
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 10894 117854 18064
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 17940
rect 122606 17509 122666 19350
rect 124674 18023 125294 18064
rect 124674 17787 124706 18023
rect 124942 17787 125026 18023
rect 125262 17787 125294 18023
rect 125918 17917 125978 19350
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 125915 17916 125981 17917
rect 125915 17852 125916 17916
rect 125980 17852 125981 17916
rect 125915 17851 125981 17852
rect 122603 17508 122669 17509
rect 122603 17444 122604 17508
rect 122668 17444 122669 17508
rect 122603 17443 122669 17444
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 -4186 125294 17787
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 145794 3454 146414 18064
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 7174 150134 18064
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 10894 153854 18064
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 18064
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 164394 598054 165014 633498
rect 164394 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 165014 598054
rect 164394 597734 165014 597818
rect 164394 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 165014 597734
rect 164394 562054 165014 597498
rect 164394 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 165014 562054
rect 164394 561734 165014 561818
rect 164394 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 165014 561734
rect 164394 526054 165014 561498
rect 164394 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 165014 526054
rect 164394 525734 165014 525818
rect 164394 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 165014 525734
rect 164394 490054 165014 525498
rect 164394 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 165014 490054
rect 164394 489734 165014 489818
rect 164394 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 165014 489734
rect 164394 454054 165014 489498
rect 164394 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 165014 454054
rect 164394 453734 165014 453818
rect 164394 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 165014 453734
rect 164394 418054 165014 453498
rect 164394 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 165014 418054
rect 164394 417734 165014 417818
rect 164394 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 165014 417734
rect 164394 382054 165014 417498
rect 164394 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 165014 382054
rect 164394 381734 165014 381818
rect 164394 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 165014 381734
rect 164394 346054 165014 381498
rect 164394 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 165014 346054
rect 164394 345734 165014 345818
rect 164394 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 165014 345734
rect 164394 310054 165014 345498
rect 164394 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 165014 310054
rect 164394 309734 165014 309818
rect 164394 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 165014 309734
rect 164394 274054 165014 309498
rect 164394 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 165014 274054
rect 164394 273734 165014 273818
rect 164394 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 165014 273734
rect 164394 238054 165014 273498
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 130054 165014 165498
rect 164394 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 165014 130054
rect 164394 129734 165014 129818
rect 164394 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 165014 129734
rect 164394 94054 165014 129498
rect 164394 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 165014 94054
rect 164394 93734 165014 93818
rect 164394 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 165014 93734
rect 164394 58054 165014 93498
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 168114 601774 168734 637218
rect 168114 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 168734 601774
rect 168114 601454 168734 601538
rect 168114 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 168734 601454
rect 168114 565774 168734 601218
rect 168114 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 168734 565774
rect 168114 565454 168734 565538
rect 168114 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 168734 565454
rect 168114 529774 168734 565218
rect 168114 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 168734 529774
rect 168114 529454 168734 529538
rect 168114 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 168734 529454
rect 168114 493774 168734 529218
rect 168114 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 168734 493774
rect 168114 493454 168734 493538
rect 168114 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 168734 493454
rect 168114 457774 168734 493218
rect 168114 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 168734 457774
rect 168114 457454 168734 457538
rect 168114 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 168734 457454
rect 168114 421774 168734 457218
rect 168114 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 168734 421774
rect 168114 421454 168734 421538
rect 168114 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 168734 421454
rect 168114 385774 168734 421218
rect 168114 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 168734 385774
rect 168114 385454 168734 385538
rect 168114 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 168734 385454
rect 168114 349774 168734 385218
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 168114 313774 168734 349218
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 168114 277774 168734 313218
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 168114 241774 168734 277218
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 168114 205774 168734 241218
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 168114 169774 168734 205218
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 97774 168734 133218
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 168114 61774 168734 97218
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 168114 25774 168734 61218
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 641494 172454 676938
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 605494 172454 640938
rect 171834 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 172454 605494
rect 171834 605174 172454 605258
rect 171834 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 172454 605174
rect 171834 569494 172454 604938
rect 171834 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 172454 569494
rect 171834 569174 172454 569258
rect 171834 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 172454 569174
rect 171834 533494 172454 568938
rect 171834 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 172454 533494
rect 171834 533174 172454 533258
rect 171834 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 172454 533174
rect 171834 497494 172454 532938
rect 171834 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 172454 497494
rect 171834 497174 172454 497258
rect 171834 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 172454 497174
rect 171834 461494 172454 496938
rect 171834 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 172454 461494
rect 171834 461174 172454 461258
rect 171834 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 172454 461174
rect 171834 425494 172454 460938
rect 171834 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 172454 425494
rect 171834 425174 172454 425258
rect 171834 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 172454 425174
rect 171834 389494 172454 424938
rect 171834 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 172454 389494
rect 171834 389174 172454 389258
rect 171834 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 172454 389174
rect 171834 353494 172454 388938
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 171834 317494 172454 352938
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 171834 281494 172454 316938
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 171834 245494 172454 280938
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 171834 209494 172454 244938
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 171834 173494 172454 208938
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 171834 101494 172454 136938
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 171834 65494 172454 100938
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 171834 29494 172454 64938
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 184059 457196 184125 457197
rect 184059 457132 184060 457196
rect 184124 457132 184125 457196
rect 184059 457131 184125 457132
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 184062 106861 184122 457131
rect 184243 455836 184309 455837
rect 184243 455772 184244 455836
rect 184308 455772 184309 455836
rect 184243 455771 184309 455772
rect 184246 108493 184306 455771
rect 185163 453252 185229 453253
rect 185163 453188 185164 453252
rect 185228 453188 185229 453252
rect 185163 453187 185229 453188
rect 184243 108492 184309 108493
rect 184243 108428 184244 108492
rect 184308 108428 184309 108492
rect 184243 108427 184309 108428
rect 184059 106860 184125 106861
rect 184059 106796 184060 106860
rect 184124 106796 184125 106860
rect 184059 106795 184125 106796
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 185166 19277 185226 453187
rect 185514 439174 186134 474618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 188475 458964 188541 458965
rect 188475 458900 188476 458964
rect 188540 458900 188541 458964
rect 188475 458899 188541 458900
rect 186819 457332 186885 457333
rect 186819 457268 186820 457332
rect 186884 457268 186885 457332
rect 186819 457267 186885 457268
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 186822 108765 186882 457267
rect 187003 456108 187069 456109
rect 187003 456044 187004 456108
rect 187068 456044 187069 456108
rect 187003 456043 187069 456044
rect 186819 108764 186885 108765
rect 186819 108700 186820 108764
rect 186884 108700 186885 108764
rect 186819 108699 186885 108700
rect 187006 107133 187066 456043
rect 187187 455972 187253 455973
rect 187187 455908 187188 455972
rect 187252 455908 187253 455972
rect 187187 455907 187253 455908
rect 187190 108629 187250 455907
rect 188291 454612 188357 454613
rect 188291 454548 188292 454612
rect 188356 454548 188357 454612
rect 188291 454547 188357 454548
rect 187371 450396 187437 450397
rect 187371 450332 187372 450396
rect 187436 450332 187437 450396
rect 187371 450331 187437 450332
rect 187187 108628 187253 108629
rect 187187 108564 187188 108628
rect 187252 108564 187253 108628
rect 187187 108563 187253 108564
rect 187374 107269 187434 450331
rect 187371 107268 187437 107269
rect 187371 107204 187372 107268
rect 187436 107204 187437 107268
rect 187371 107203 187437 107204
rect 187003 107132 187069 107133
rect 187003 107068 187004 107132
rect 187068 107068 187069 107132
rect 187003 107067 187069 107068
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185163 19276 185229 19277
rect 185163 19212 185164 19276
rect 185228 19212 185229 19276
rect 185163 19211 185229 19212
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 7174 186134 42618
rect 188294 17645 188354 454547
rect 188478 108901 188538 458899
rect 188843 451484 188909 451485
rect 188843 451420 188844 451484
rect 188908 451420 188909 451484
rect 188843 451419 188909 451420
rect 188659 451348 188725 451349
rect 188659 451284 188660 451348
rect 188724 451284 188725 451348
rect 188659 451283 188725 451284
rect 188475 108900 188541 108901
rect 188475 108836 188476 108900
rect 188540 108836 188541 108900
rect 188475 108835 188541 108836
rect 188662 105501 188722 451283
rect 188846 105637 188906 451419
rect 189234 442894 189854 478338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 195835 680372 195901 680373
rect 195835 680308 195836 680372
rect 195900 680308 195901 680372
rect 195835 680307 195901 680308
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 195099 587348 195165 587349
rect 195099 587284 195100 587348
rect 195164 587284 195165 587348
rect 195099 587283 195165 587284
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192707 463724 192773 463725
rect 192707 463660 192708 463724
rect 192772 463660 192773 463724
rect 192707 463659 192773 463660
rect 192155 461412 192221 461413
rect 192155 461348 192156 461412
rect 192220 461348 192221 461412
rect 192155 461347 192221 461348
rect 190315 454748 190381 454749
rect 190315 454684 190316 454748
rect 190380 454684 190381 454748
rect 190315 454683 190381 454684
rect 190131 449716 190197 449717
rect 190131 449652 190132 449716
rect 190196 449652 190197 449716
rect 190131 449651 190197 449652
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 190134 249117 190194 449651
rect 190131 249116 190197 249117
rect 190131 249052 190132 249116
rect 190196 249052 190197 249116
rect 190131 249051 190197 249052
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 188843 105636 188909 105637
rect 188843 105572 188844 105636
rect 188908 105572 188909 105636
rect 188843 105571 188909 105572
rect 188659 105500 188725 105501
rect 188659 105436 188660 105500
rect 188724 105436 188725 105500
rect 188659 105435 188725 105436
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 188291 17644 188357 17645
rect 188291 17580 188292 17644
rect 188356 17580 188357 17644
rect 188291 17579 188357 17580
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 10894 189854 46338
rect 190318 30021 190378 454683
rect 191051 454476 191117 454477
rect 191051 454412 191052 454476
rect 191116 454412 191117 454476
rect 191051 454411 191117 454412
rect 190315 30020 190381 30021
rect 190315 29956 190316 30020
rect 190380 29956 190381 30020
rect 190315 29955 190381 29956
rect 191054 17509 191114 454411
rect 191603 451348 191669 451349
rect 191603 451284 191604 451348
rect 191668 451284 191669 451348
rect 191603 451283 191669 451284
rect 191235 450804 191301 450805
rect 191235 450740 191236 450804
rect 191300 450740 191301 450804
rect 191235 450739 191301 450740
rect 191238 107405 191298 450739
rect 191419 450532 191485 450533
rect 191419 450468 191420 450532
rect 191484 450468 191485 450532
rect 191419 450467 191485 450468
rect 191235 107404 191301 107405
rect 191235 107340 191236 107404
rect 191300 107340 191301 107404
rect 191235 107339 191301 107340
rect 191422 106997 191482 450467
rect 191419 106996 191485 106997
rect 191419 106932 191420 106996
rect 191484 106932 191485 106996
rect 191419 106931 191485 106932
rect 191606 105773 191666 451283
rect 192158 369885 192218 461347
rect 192523 453116 192589 453117
rect 192523 453052 192524 453116
rect 192588 453052 192589 453116
rect 192523 453051 192589 453052
rect 192339 450668 192405 450669
rect 192339 450604 192340 450668
rect 192404 450604 192405 450668
rect 192339 450603 192405 450604
rect 192342 395997 192402 450603
rect 192339 395996 192405 395997
rect 192339 395932 192340 395996
rect 192404 395932 192405 395996
rect 192339 395931 192405 395932
rect 192339 394772 192405 394773
rect 192339 394708 192340 394772
rect 192404 394708 192405 394772
rect 192339 394707 192405 394708
rect 192155 369884 192221 369885
rect 192155 369820 192156 369884
rect 192220 369820 192221 369884
rect 192155 369819 192221 369820
rect 191787 369204 191853 369205
rect 191787 369140 191788 369204
rect 191852 369140 191853 369204
rect 191787 369139 191853 369140
rect 191603 105772 191669 105773
rect 191603 105708 191604 105772
rect 191668 105708 191669 105772
rect 191603 105707 191669 105708
rect 191051 17508 191117 17509
rect 191051 17444 191052 17508
rect 191116 17444 191117 17508
rect 191051 17443 191117 17444
rect 191790 17101 191850 369139
rect 192342 17781 192402 394707
rect 192339 17780 192405 17781
rect 192339 17716 192340 17780
rect 192404 17716 192405 17780
rect 192339 17715 192405 17716
rect 192526 17645 192586 453051
rect 192523 17644 192589 17645
rect 192523 17580 192524 17644
rect 192588 17580 192589 17644
rect 192523 17579 192589 17580
rect 192710 17237 192770 463659
rect 192954 446614 193574 482058
rect 195102 475421 195162 587283
rect 195838 497997 195898 680307
rect 196674 666334 197294 708122
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 199331 700364 199397 700365
rect 199331 700300 199332 700364
rect 199396 700300 199397 700364
rect 199331 700299 199397 700300
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 630334 197294 665778
rect 196674 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 197294 630334
rect 196674 630014 197294 630098
rect 196674 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 197294 630014
rect 196674 594334 197294 629778
rect 196674 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 197294 594334
rect 196674 594014 197294 594098
rect 196674 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 197294 594014
rect 196674 558334 197294 593778
rect 198043 587212 198109 587213
rect 198043 587148 198044 587212
rect 198108 587148 198109 587212
rect 198043 587147 198109 587148
rect 197859 584628 197925 584629
rect 197859 584564 197860 584628
rect 197924 584564 197925 584628
rect 197859 584563 197925 584564
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 196674 522334 197294 557778
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 195835 497996 195901 497997
rect 195835 497932 195836 497996
rect 195900 497932 195901 497996
rect 195835 497931 195901 497932
rect 196674 486334 197294 521778
rect 196674 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 197294 486334
rect 196674 486014 197294 486098
rect 196674 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 197294 486014
rect 195099 475420 195165 475421
rect 195099 475356 195100 475420
rect 195164 475356 195165 475420
rect 195099 475355 195165 475356
rect 196674 450334 197294 485778
rect 197862 460189 197922 584563
rect 198046 465901 198106 587147
rect 199334 468485 199394 700299
rect 199883 680508 199949 680509
rect 199883 680444 199884 680508
rect 199948 680444 199949 680508
rect 199883 680443 199949 680444
rect 199515 585716 199581 585717
rect 199515 585652 199516 585716
rect 199580 585652 199581 585716
rect 199515 585651 199581 585652
rect 199518 499493 199578 585651
rect 199699 584356 199765 584357
rect 199699 584292 199700 584356
rect 199764 584292 199765 584356
rect 199699 584291 199765 584292
rect 199702 577010 199762 584291
rect 199886 577149 199946 680443
rect 200394 670054 201014 709082
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 203195 700908 203261 700909
rect 203195 700844 203196 700908
rect 203260 700844 203261 700908
rect 203195 700843 203261 700844
rect 202459 700772 202525 700773
rect 202459 700708 202460 700772
rect 202524 700708 202525 700772
rect 202459 700707 202525 700708
rect 202275 700636 202341 700637
rect 202275 700572 202276 700636
rect 202340 700572 202341 700636
rect 202275 700571 202341 700572
rect 202091 700500 202157 700501
rect 202091 700436 202092 700500
rect 202156 700436 202157 700500
rect 202091 700435 202157 700436
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 598054 201014 633498
rect 200394 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 201014 598054
rect 200394 597734 201014 597818
rect 200394 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 201014 597734
rect 199883 577148 199949 577149
rect 199883 577084 199884 577148
rect 199948 577084 199949 577148
rect 199883 577083 199949 577084
rect 199702 576950 200130 577010
rect 199883 576876 199949 576877
rect 199883 576870 199884 576876
rect 199702 576812 199884 576870
rect 199948 576812 199949 576876
rect 199702 576811 199949 576812
rect 199702 576810 199946 576811
rect 199702 509690 199762 576810
rect 200070 576330 200130 576950
rect 199886 576270 200130 576330
rect 199886 567210 199946 576270
rect 199886 567150 200130 567210
rect 200070 566810 200130 567150
rect 199886 566750 200130 566810
rect 199886 557970 199946 566750
rect 200394 562054 201014 597498
rect 201355 584492 201421 584493
rect 201355 584428 201356 584492
rect 201420 584428 201421 584492
rect 201355 584427 201421 584428
rect 200394 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 201014 562054
rect 200394 561734 201014 561818
rect 200394 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 201014 561734
rect 199886 557910 200130 557970
rect 200070 557550 200130 557910
rect 199886 557490 200130 557550
rect 199886 547890 199946 557490
rect 199886 547830 200130 547890
rect 200070 547770 200130 547830
rect 199886 547710 200130 547770
rect 199886 538930 199946 547710
rect 199886 538870 200314 538930
rect 200254 538230 200314 538870
rect 199886 538170 200314 538230
rect 199886 528570 199946 538170
rect 199886 528510 200130 528570
rect 200070 528050 200130 528510
rect 199886 527990 200130 528050
rect 199886 519210 199946 527990
rect 200394 526054 201014 561498
rect 200394 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 201014 526054
rect 200394 525734 201014 525818
rect 200394 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 201014 525734
rect 199886 519150 200130 519210
rect 200070 518910 200130 519150
rect 199886 518850 200130 518910
rect 199886 514770 199946 518850
rect 199886 514710 200130 514770
rect 199702 509630 199946 509690
rect 199699 505204 199765 505205
rect 199699 505140 199700 505204
rect 199764 505140 199765 505204
rect 199699 505139 199765 505140
rect 199702 499629 199762 505139
rect 199699 499628 199765 499629
rect 199699 499564 199700 499628
rect 199764 499564 199765 499628
rect 199699 499563 199765 499564
rect 199515 499492 199581 499493
rect 199515 499428 199516 499492
rect 199580 499428 199581 499492
rect 199515 499427 199581 499428
rect 199886 497861 199946 509630
rect 200070 505205 200130 514710
rect 200067 505204 200133 505205
rect 200067 505140 200068 505204
rect 200132 505140 200133 505204
rect 200067 505139 200133 505140
rect 200067 499628 200133 499629
rect 200067 499564 200068 499628
rect 200132 499590 200133 499628
rect 200132 499564 200314 499590
rect 200067 499563 200314 499564
rect 200070 499530 200314 499563
rect 199883 497860 199949 497861
rect 199883 497796 199884 497860
rect 199948 497796 199949 497860
rect 199883 497795 199949 497796
rect 200254 497450 200314 499530
rect 199886 497390 200314 497450
rect 199331 468484 199397 468485
rect 199331 468420 199332 468484
rect 199396 468420 199397 468484
rect 199331 468419 199397 468420
rect 198043 465900 198109 465901
rect 198043 465836 198044 465900
rect 198108 465836 198109 465900
rect 198043 465835 198109 465836
rect 199886 461685 199946 497390
rect 200394 490054 201014 525498
rect 200394 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 201014 490054
rect 200394 489734 201014 489818
rect 200394 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 201014 489734
rect 199883 461684 199949 461685
rect 199883 461620 199884 461684
rect 199948 461620 199949 461684
rect 199883 461619 199949 461620
rect 197859 460188 197925 460189
rect 197859 460124 197860 460188
rect 197924 460124 197925 460188
rect 197859 460123 197925 460124
rect 193811 450260 193877 450261
rect 193811 450196 193812 450260
rect 193876 450196 193877 450260
rect 193811 450195 193877 450196
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 193814 193901 193874 450195
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 193995 449308 194061 449309
rect 193995 449244 193996 449308
rect 194060 449244 194061 449308
rect 193995 449243 194061 449244
rect 193998 194037 194058 449243
rect 194208 435454 194528 435486
rect 194208 435218 194250 435454
rect 194486 435218 194528 435454
rect 194208 435134 194528 435218
rect 194208 434898 194250 435134
rect 194486 434898 194528 435134
rect 194208 434866 194528 434898
rect 196674 414334 197294 449778
rect 196674 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 197294 414334
rect 196674 414014 197294 414098
rect 196674 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 197294 414014
rect 194208 399454 194528 399486
rect 194208 399218 194250 399454
rect 194486 399218 194528 399454
rect 194208 399134 194528 399218
rect 194208 398898 194250 399134
rect 194486 398898 194528 399134
rect 194208 398866 194528 398898
rect 196674 378334 197294 413778
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 194208 363454 194528 363486
rect 194208 363218 194250 363454
rect 194486 363218 194528 363454
rect 194208 363134 194528 363218
rect 194208 362898 194250 363134
rect 194486 362898 194528 363134
rect 194208 362866 194528 362898
rect 196674 342334 197294 377778
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 194208 327454 194528 327486
rect 194208 327218 194250 327454
rect 194486 327218 194528 327454
rect 194208 327134 194528 327218
rect 194208 326898 194250 327134
rect 194486 326898 194528 327134
rect 194208 326866 194528 326898
rect 196674 306334 197294 341778
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 194208 291454 194528 291486
rect 194208 291218 194250 291454
rect 194486 291218 194528 291454
rect 194208 291134 194528 291218
rect 194208 290898 194250 291134
rect 194486 290898 194528 291134
rect 194208 290866 194528 290898
rect 196674 270334 197294 305778
rect 196674 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 197294 270334
rect 196674 270014 197294 270098
rect 196674 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 197294 270014
rect 194208 255454 194528 255486
rect 194208 255218 194250 255454
rect 194486 255218 194528 255454
rect 194208 255134 194528 255218
rect 194208 254898 194250 255134
rect 194486 254898 194528 255134
rect 194208 254866 194528 254898
rect 196674 234334 197294 269778
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 196674 198334 197294 233778
rect 196674 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 197294 198334
rect 196674 198014 197294 198098
rect 196674 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 197294 198014
rect 193995 194036 194061 194037
rect 193995 193972 193996 194036
rect 194060 193972 194061 194036
rect 193995 193971 194061 193972
rect 193811 193900 193877 193901
rect 193811 193836 193812 193900
rect 193876 193836 193877 193900
rect 193811 193835 193877 193836
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192707 17236 192773 17237
rect 192707 17172 192708 17236
rect 192772 17172 192773 17236
rect 192707 17171 192773 17172
rect 191787 17100 191853 17101
rect 191787 17036 191788 17100
rect 191852 17036 191853 17100
rect 191787 17035 191853 17036
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 162334 197294 197778
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 196674 126334 197294 161778
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 196674 90334 197294 125778
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 196674 54334 197294 89778
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 454054 201014 489498
rect 201358 461549 201418 584427
rect 202094 500581 202154 700435
rect 202278 500717 202338 700571
rect 202462 500853 202522 700707
rect 202643 700364 202709 700365
rect 202643 700300 202644 700364
rect 202708 700300 202709 700364
rect 202643 700299 202709 700300
rect 202459 500852 202525 500853
rect 202459 500788 202460 500852
rect 202524 500788 202525 500852
rect 202459 500787 202525 500788
rect 202275 500716 202341 500717
rect 202275 500652 202276 500716
rect 202340 500652 202341 500716
rect 202275 500651 202341 500652
rect 202091 500580 202157 500581
rect 202091 500516 202092 500580
rect 202156 500516 202157 500580
rect 202091 500515 202157 500516
rect 202646 499901 202706 700299
rect 203198 500037 203258 700843
rect 203563 682684 203629 682685
rect 203563 682620 203564 682684
rect 203628 682620 203629 682684
rect 203563 682619 203629 682620
rect 203379 682412 203445 682413
rect 203379 682348 203380 682412
rect 203444 682348 203445 682412
rect 203379 682347 203445 682348
rect 203382 500445 203442 682347
rect 203379 500444 203445 500445
rect 203379 500380 203380 500444
rect 203444 500380 203445 500444
rect 203379 500379 203445 500380
rect 203195 500036 203261 500037
rect 203195 499972 203196 500036
rect 203260 499972 203261 500036
rect 203195 499971 203261 499972
rect 202643 499900 202709 499901
rect 202643 499836 202644 499900
rect 202708 499836 202709 499900
rect 202643 499835 202709 499836
rect 203566 466173 203626 682619
rect 203747 682548 203813 682549
rect 203747 682484 203748 682548
rect 203812 682484 203813 682548
rect 203747 682483 203813 682484
rect 203563 466172 203629 466173
rect 203563 466108 203564 466172
rect 203628 466108 203629 466172
rect 203563 466107 203629 466108
rect 201355 461548 201421 461549
rect 201355 461484 201356 461548
rect 201420 461484 201421 461548
rect 201355 461483 201421 461484
rect 200394 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 201014 454054
rect 200394 453734 201014 453818
rect 200394 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 201014 453734
rect 200394 418054 201014 453498
rect 203750 452165 203810 682483
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 204208 651454 204528 651486
rect 204208 651218 204250 651454
rect 204486 651218 204528 651454
rect 204208 651134 204528 651218
rect 204208 650898 204250 651134
rect 204486 650898 204528 651134
rect 204208 650866 204528 650898
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 204208 615454 204528 615486
rect 204208 615218 204250 615454
rect 204486 615218 204528 615454
rect 204208 615134 204528 615218
rect 204208 614898 204250 615134
rect 204486 614898 204528 615134
rect 204208 614866 204528 614898
rect 207834 605494 208454 640938
rect 207834 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 208454 605494
rect 207834 605174 208454 605258
rect 207834 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 208454 605174
rect 204208 579454 204528 579486
rect 204208 579218 204250 579454
rect 204486 579218 204528 579454
rect 204208 579134 204528 579218
rect 204208 578898 204250 579134
rect 204486 578898 204528 579134
rect 204208 578866 204528 578898
rect 207834 569494 208454 604938
rect 207834 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 208454 569494
rect 207834 569174 208454 569258
rect 207834 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 208454 569174
rect 204208 543454 204528 543486
rect 204208 543218 204250 543454
rect 204486 543218 204528 543454
rect 204208 543134 204528 543218
rect 204208 542898 204250 543134
rect 204486 542898 204528 543134
rect 204208 542866 204528 542898
rect 207834 533494 208454 568938
rect 207834 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 208454 533494
rect 207834 533174 208454 533258
rect 207834 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 208454 533174
rect 204208 507454 204528 507486
rect 204208 507218 204250 507454
rect 204486 507218 204528 507454
rect 204208 507134 204528 507218
rect 204208 506898 204250 507134
rect 204486 506898 204528 507134
rect 204208 506866 204528 506898
rect 204114 493774 204734 500068
rect 204114 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 204734 493774
rect 204114 493454 204734 493538
rect 204114 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 204734 493454
rect 204114 457774 204734 493218
rect 204114 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 204734 457774
rect 204114 457454 204734 457538
rect 204114 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 204734 457454
rect 203747 452164 203813 452165
rect 203747 452100 203748 452164
rect 203812 452100 203813 452164
rect 203747 452099 203813 452100
rect 200394 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 201014 418054
rect 200394 417734 201014 417818
rect 200394 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 201014 417734
rect 200394 382054 201014 417498
rect 200394 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 201014 382054
rect 200394 381734 201014 381818
rect 200394 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 201014 381734
rect 200394 346054 201014 381498
rect 200394 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 201014 346054
rect 200394 345734 201014 345818
rect 200394 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 201014 345734
rect 200394 310054 201014 345498
rect 200394 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 201014 310054
rect 200394 309734 201014 309818
rect 200394 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 201014 309734
rect 200394 274054 201014 309498
rect 200394 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 201014 274054
rect 200394 273734 201014 273818
rect 200394 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 201014 273734
rect 200394 238054 201014 273498
rect 200394 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 201014 238054
rect 200394 237734 201014 237818
rect 200394 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 201014 237734
rect 200394 202054 201014 237498
rect 200394 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 201014 202054
rect 200394 201734 201014 201818
rect 200394 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 201014 201734
rect 200394 166054 201014 201498
rect 200394 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 201014 166054
rect 200394 165734 201014 165818
rect 200394 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 201014 165734
rect 200394 130054 201014 165498
rect 200394 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 201014 130054
rect 200394 129734 201014 129818
rect 200394 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 201014 129734
rect 200394 94054 201014 129498
rect 200394 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 201014 94054
rect 200394 93734 201014 93818
rect 200394 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 201014 93734
rect 200394 58054 201014 93498
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 421774 204734 457218
rect 204114 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 204734 421774
rect 204114 421454 204734 421538
rect 204114 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 204734 421454
rect 204114 385774 204734 421218
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 204114 349774 204734 385218
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 204114 313774 204734 349218
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 204114 277774 204734 313218
rect 204114 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 204734 277774
rect 204114 277454 204734 277538
rect 204114 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 204734 277454
rect 204114 241774 204734 277218
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 204114 205774 204734 241218
rect 204114 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 204734 205774
rect 204114 205454 204734 205538
rect 204114 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 204734 205454
rect 204114 169774 204734 205218
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 204114 133774 204734 169218
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 204114 97774 204734 133218
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 204114 61774 204734 97218
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 204114 25774 204734 61218
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 497494 208454 532938
rect 207834 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 208454 497494
rect 207834 497174 208454 497258
rect 207834 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 208454 497174
rect 207834 461494 208454 496938
rect 207834 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 208454 461494
rect 207834 461174 208454 461258
rect 207834 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 208454 461174
rect 207834 425494 208454 460938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 219568 655174 219888 655206
rect 219568 654938 219610 655174
rect 219846 654938 219888 655174
rect 219568 654854 219888 654938
rect 219568 654618 219610 654854
rect 219846 654618 219888 654854
rect 219568 654586 219888 654618
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 219568 619174 219888 619206
rect 219568 618938 219610 619174
rect 219846 618938 219888 619174
rect 219568 618854 219888 618938
rect 219568 618618 219610 618854
rect 219846 618618 219888 618854
rect 219568 618586 219888 618618
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 219568 583174 219888 583206
rect 219568 582938 219610 583174
rect 219846 582938 219888 583174
rect 219568 582854 219888 582938
rect 219568 582618 219610 582854
rect 219846 582618 219888 582854
rect 219568 582586 219888 582618
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 219568 547174 219888 547206
rect 219568 546938 219610 547174
rect 219846 546938 219888 547174
rect 219568 546854 219888 546938
rect 219568 546618 219610 546854
rect 219846 546618 219888 546854
rect 219568 546586 219888 546618
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 219568 511174 219888 511206
rect 219568 510938 219610 511174
rect 219846 510938 219888 511174
rect 219568 510854 219888 510938
rect 219568 510618 219610 510854
rect 219846 510618 219888 510854
rect 219568 510586 219888 510618
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 209568 439174 209888 439206
rect 209568 438938 209610 439174
rect 209846 438938 209888 439174
rect 209568 438854 209888 438938
rect 209568 438618 209610 438854
rect 209846 438618 209888 438854
rect 209568 438586 209888 438618
rect 207834 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 208454 425494
rect 207834 425174 208454 425258
rect 207834 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 208454 425174
rect 207834 389494 208454 424938
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 209568 403174 209888 403206
rect 209568 402938 209610 403174
rect 209846 402938 209888 403174
rect 209568 402854 209888 402938
rect 209568 402618 209610 402854
rect 209846 402618 209888 402854
rect 209568 402586 209888 402618
rect 207834 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 208454 389494
rect 207834 389174 208454 389258
rect 207834 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 208454 389174
rect 207834 353494 208454 388938
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 209568 367174 209888 367206
rect 209568 366938 209610 367174
rect 209846 366938 209888 367174
rect 209568 366854 209888 366938
rect 209568 366618 209610 366854
rect 209846 366618 209888 366854
rect 209568 366586 209888 366618
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 207834 317494 208454 352938
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 209568 331174 209888 331206
rect 209568 330938 209610 331174
rect 209846 330938 209888 331174
rect 209568 330854 209888 330938
rect 209568 330618 209610 330854
rect 209846 330618 209888 330854
rect 209568 330586 209888 330618
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 207834 281494 208454 316938
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 209568 295174 209888 295206
rect 209568 294938 209610 295174
rect 209846 294938 209888 295174
rect 209568 294854 209888 294938
rect 209568 294618 209610 294854
rect 209846 294618 209888 294854
rect 209568 294586 209888 294618
rect 207834 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 208454 281494
rect 207834 281174 208454 281258
rect 207834 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 208454 281174
rect 207834 245494 208454 280938
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 209568 259174 209888 259206
rect 209568 258938 209610 259174
rect 209846 258938 209888 259174
rect 209568 258854 209888 258938
rect 209568 258618 209610 258854
rect 209846 258618 209888 258854
rect 209568 258586 209888 258618
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 207834 209494 208454 244938
rect 207834 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 208454 209494
rect 207834 209174 208454 209258
rect 207834 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 208454 209174
rect 207834 173494 208454 208938
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 207834 137494 208454 172938
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 207834 101494 208454 136938
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 105244 218414 110898
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 449580 225854 478338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 224928 435454 225248 435486
rect 224928 435218 224970 435454
rect 225206 435218 225248 435454
rect 224928 435134 225248 435218
rect 224928 434898 224970 435134
rect 225206 434898 225248 435134
rect 224928 434866 225248 434898
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 224928 399454 225248 399486
rect 224928 399218 224970 399454
rect 225206 399218 225248 399454
rect 224928 399134 225248 399218
rect 224928 398898 224970 399134
rect 225206 398898 225248 399134
rect 224928 398866 225248 398898
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 224928 363454 225248 363486
rect 224928 363218 224970 363454
rect 225206 363218 225248 363454
rect 224928 363134 225248 363218
rect 224928 362898 224970 363134
rect 225206 362898 225248 363134
rect 224928 362866 225248 362898
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 224928 327454 225248 327486
rect 224928 327218 224970 327454
rect 225206 327218 225248 327454
rect 224928 327134 225248 327218
rect 224928 326898 224970 327134
rect 225206 326898 225248 327134
rect 224928 326866 225248 326898
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 224928 291454 225248 291486
rect 224928 291218 224970 291454
rect 225206 291218 225248 291454
rect 224928 291134 225248 291218
rect 224928 290898 224970 291134
rect 225206 290898 225248 291134
rect 224928 290866 225248 290898
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 224928 255454 225248 255486
rect 224928 255218 224970 255454
rect 225206 255218 225248 255454
rect 224928 255134 225248 255218
rect 224928 254898 224970 255134
rect 225206 254898 225248 255134
rect 224928 254866 225248 254898
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 105244 222134 114618
rect 225234 226894 225854 250068
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 105244 225854 118338
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 105244 229574 122058
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 630334 233294 665778
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 234928 651454 235248 651486
rect 234928 651218 234970 651454
rect 235206 651218 235248 651454
rect 234928 651134 235248 651218
rect 234928 650898 234970 651134
rect 235206 650898 235248 651134
rect 234928 650866 235248 650898
rect 232674 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 233294 630334
rect 232674 630014 233294 630098
rect 232674 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 233294 630014
rect 232674 594334 233294 629778
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 234928 615454 235248 615486
rect 234928 615218 234970 615454
rect 235206 615218 235248 615454
rect 234928 615134 235248 615218
rect 234928 614898 234970 615134
rect 235206 614898 235248 615134
rect 234928 614866 235248 614898
rect 232674 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 233294 594334
rect 232674 594014 233294 594098
rect 232674 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 233294 594014
rect 232674 558334 233294 593778
rect 236394 598054 237014 633498
rect 236394 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 237014 598054
rect 236394 597734 237014 597818
rect 236394 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 237014 597734
rect 234928 579454 235248 579486
rect 234928 579218 234970 579454
rect 235206 579218 235248 579454
rect 234928 579134 235248 579218
rect 234928 578898 234970 579134
rect 235206 578898 235248 579134
rect 234928 578866 235248 578898
rect 232674 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 233294 558334
rect 232674 558014 233294 558098
rect 232674 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 233294 558014
rect 232674 522334 233294 557778
rect 236394 562054 237014 597498
rect 236394 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 237014 562054
rect 236394 561734 237014 561818
rect 236394 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 237014 561734
rect 234928 543454 235248 543486
rect 234928 543218 234970 543454
rect 235206 543218 235248 543454
rect 234928 543134 235248 543218
rect 234928 542898 234970 543134
rect 235206 542898 235248 543134
rect 234928 542866 235248 542898
rect 232674 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 233294 522334
rect 232674 522014 233294 522098
rect 232674 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 233294 522014
rect 232674 486334 233294 521778
rect 236394 526054 237014 561498
rect 236394 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 237014 526054
rect 236394 525734 237014 525818
rect 236394 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 237014 525734
rect 234928 507454 235248 507486
rect 234928 507218 234970 507454
rect 235206 507218 235248 507454
rect 234928 507134 235248 507218
rect 234928 506898 234970 507134
rect 235206 506898 235248 507134
rect 234928 506866 235248 506898
rect 232674 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 233294 486334
rect 232674 486014 233294 486098
rect 232674 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 233294 486014
rect 232674 450334 233294 485778
rect 232674 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 233294 450334
rect 232674 450014 233294 450098
rect 232674 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 233294 450014
rect 232674 414334 233294 449778
rect 232674 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 233294 414334
rect 232674 414014 233294 414098
rect 232674 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 233294 414014
rect 232674 378334 233294 413778
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 232674 342334 233294 377778
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 232674 306334 233294 341778
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 232674 270334 233294 305778
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 232674 234334 233294 269778
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 232674 198334 233294 233778
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 232674 162334 233294 197778
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 232674 126334 233294 161778
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 232674 105244 233294 125778
rect 236394 490054 237014 525498
rect 236394 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 237014 490054
rect 236394 489734 237014 489818
rect 236394 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 237014 489734
rect 236394 454054 237014 489498
rect 236394 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 237014 454054
rect 236394 453734 237014 453818
rect 236394 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 237014 453734
rect 236394 418054 237014 453498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 678961 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 678961 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 678961 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264467 679692 264533 679693
rect 264467 679628 264468 679692
rect 264532 679628 264533 679692
rect 264467 679627 264533 679628
rect 264470 678333 264530 679627
rect 264954 678961 265574 698058
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 269251 679692 269317 679693
rect 269251 679628 269252 679692
rect 269316 679628 269317 679692
rect 269251 679627 269317 679628
rect 264467 678332 264533 678333
rect 264467 678268 264468 678332
rect 264532 678268 264533 678332
rect 264467 678267 264533 678268
rect 269254 678197 269314 679627
rect 289794 678961 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 678961 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 678961 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 678961 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 678961 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 678961 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 269251 678196 269317 678197
rect 269251 678132 269252 678196
rect 269316 678132 269317 678196
rect 269251 678131 269317 678132
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 250288 655174 250608 655206
rect 250288 654938 250330 655174
rect 250566 654938 250608 655174
rect 250288 654854 250608 654938
rect 250288 654618 250330 654854
rect 250566 654618 250608 654854
rect 250288 654586 250608 654618
rect 281008 655174 281328 655206
rect 281008 654938 281050 655174
rect 281286 654938 281328 655174
rect 281008 654854 281328 654938
rect 281008 654618 281050 654854
rect 281286 654618 281328 654854
rect 281008 654586 281328 654618
rect 311728 655174 312048 655206
rect 311728 654938 311770 655174
rect 312006 654938 312048 655174
rect 311728 654854 312048 654938
rect 311728 654618 311770 654854
rect 312006 654618 312048 654854
rect 311728 654586 312048 654618
rect 265648 651454 265968 651486
rect 265648 651218 265690 651454
rect 265926 651218 265968 651454
rect 265648 651134 265968 651218
rect 265648 650898 265690 651134
rect 265926 650898 265968 651134
rect 265648 650866 265968 650898
rect 296368 651454 296688 651486
rect 296368 651218 296410 651454
rect 296646 651218 296688 651454
rect 296368 651134 296688 651218
rect 296368 650898 296410 651134
rect 296646 650898 296688 651134
rect 296368 650866 296688 650898
rect 327088 651454 327408 651486
rect 327088 651218 327130 651454
rect 327366 651218 327408 651454
rect 327088 651134 327408 651218
rect 327088 650898 327130 651134
rect 327366 650898 327408 651134
rect 327088 650866 327408 650898
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 240114 601774 240734 637218
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 250288 619174 250608 619206
rect 250288 618938 250330 619174
rect 250566 618938 250608 619174
rect 250288 618854 250608 618938
rect 250288 618618 250330 618854
rect 250566 618618 250608 618854
rect 250288 618586 250608 618618
rect 281008 619174 281328 619206
rect 281008 618938 281050 619174
rect 281286 618938 281328 619174
rect 281008 618854 281328 618938
rect 281008 618618 281050 618854
rect 281286 618618 281328 618854
rect 281008 618586 281328 618618
rect 311728 619174 312048 619206
rect 311728 618938 311770 619174
rect 312006 618938 312048 619174
rect 311728 618854 312048 618938
rect 311728 618618 311770 618854
rect 312006 618618 312048 618854
rect 311728 618586 312048 618618
rect 265648 615454 265968 615486
rect 265648 615218 265690 615454
rect 265926 615218 265968 615454
rect 265648 615134 265968 615218
rect 265648 614898 265690 615134
rect 265926 614898 265968 615134
rect 265648 614866 265968 614898
rect 296368 615454 296688 615486
rect 296368 615218 296410 615454
rect 296646 615218 296688 615454
rect 296368 615134 296688 615218
rect 296368 614898 296410 615134
rect 296646 614898 296688 615134
rect 296368 614866 296688 614898
rect 327088 615454 327408 615486
rect 327088 615218 327130 615454
rect 327366 615218 327408 615454
rect 327088 615134 327408 615218
rect 327088 614898 327130 615134
rect 327366 614898 327408 615134
rect 327088 614866 327408 614898
rect 240114 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 240734 601774
rect 240114 601454 240734 601538
rect 240114 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 240734 601454
rect 240114 565774 240734 601218
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 250288 583174 250608 583206
rect 250288 582938 250330 583174
rect 250566 582938 250608 583174
rect 250288 582854 250608 582938
rect 250288 582618 250330 582854
rect 250566 582618 250608 582854
rect 250288 582586 250608 582618
rect 281008 583174 281328 583206
rect 281008 582938 281050 583174
rect 281286 582938 281328 583174
rect 281008 582854 281328 582938
rect 281008 582618 281050 582854
rect 281286 582618 281328 582854
rect 281008 582586 281328 582618
rect 311728 583174 312048 583206
rect 311728 582938 311770 583174
rect 312006 582938 312048 583174
rect 311728 582854 312048 582938
rect 311728 582618 311770 582854
rect 312006 582618 312048 582854
rect 311728 582586 312048 582618
rect 265648 579454 265968 579486
rect 265648 579218 265690 579454
rect 265926 579218 265968 579454
rect 265648 579134 265968 579218
rect 265648 578898 265690 579134
rect 265926 578898 265968 579134
rect 265648 578866 265968 578898
rect 296368 579454 296688 579486
rect 296368 579218 296410 579454
rect 296646 579218 296688 579454
rect 296368 579134 296688 579218
rect 296368 578898 296410 579134
rect 296646 578898 296688 579134
rect 296368 578866 296688 578898
rect 327088 579454 327408 579486
rect 327088 579218 327130 579454
rect 327366 579218 327408 579454
rect 327088 579134 327408 579218
rect 327088 578898 327130 579134
rect 327366 578898 327408 579134
rect 327088 578866 327408 578898
rect 240114 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 240734 565774
rect 240114 565454 240734 565538
rect 240114 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 240734 565454
rect 240114 529774 240734 565218
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 250288 547174 250608 547206
rect 250288 546938 250330 547174
rect 250566 546938 250608 547174
rect 250288 546854 250608 546938
rect 250288 546618 250330 546854
rect 250566 546618 250608 546854
rect 250288 546586 250608 546618
rect 281008 547174 281328 547206
rect 281008 546938 281050 547174
rect 281286 546938 281328 547174
rect 281008 546854 281328 546938
rect 281008 546618 281050 546854
rect 281286 546618 281328 546854
rect 281008 546586 281328 546618
rect 311728 547174 312048 547206
rect 311728 546938 311770 547174
rect 312006 546938 312048 547174
rect 311728 546854 312048 546938
rect 311728 546618 311770 546854
rect 312006 546618 312048 546854
rect 311728 546586 312048 546618
rect 265648 543454 265968 543486
rect 265648 543218 265690 543454
rect 265926 543218 265968 543454
rect 265648 543134 265968 543218
rect 265648 542898 265690 543134
rect 265926 542898 265968 543134
rect 265648 542866 265968 542898
rect 296368 543454 296688 543486
rect 296368 543218 296410 543454
rect 296646 543218 296688 543454
rect 296368 543134 296688 543218
rect 296368 542898 296410 543134
rect 296646 542898 296688 543134
rect 296368 542866 296688 542898
rect 327088 543454 327408 543486
rect 327088 543218 327130 543454
rect 327366 543218 327408 543454
rect 327088 543134 327408 543218
rect 327088 542898 327130 543134
rect 327366 542898 327408 543134
rect 327088 542866 327408 542898
rect 240114 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 240734 529774
rect 240114 529454 240734 529538
rect 240114 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 240734 529454
rect 240114 493774 240734 529218
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 250288 511174 250608 511206
rect 250288 510938 250330 511174
rect 250566 510938 250608 511174
rect 250288 510854 250608 510938
rect 250288 510618 250330 510854
rect 250566 510618 250608 510854
rect 250288 510586 250608 510618
rect 281008 511174 281328 511206
rect 281008 510938 281050 511174
rect 281286 510938 281328 511174
rect 281008 510854 281328 510938
rect 281008 510618 281050 510854
rect 281286 510618 281328 510854
rect 281008 510586 281328 510618
rect 311728 511174 312048 511206
rect 311728 510938 311770 511174
rect 312006 510938 312048 511174
rect 311728 510854 312048 510938
rect 311728 510618 311770 510854
rect 312006 510618 312048 510854
rect 311728 510586 312048 510618
rect 265648 507454 265968 507486
rect 265648 507218 265690 507454
rect 265926 507218 265968 507454
rect 265648 507134 265968 507218
rect 265648 506898 265690 507134
rect 265926 506898 265968 507134
rect 265648 506866 265968 506898
rect 296368 507454 296688 507486
rect 296368 507218 296410 507454
rect 296646 507218 296688 507454
rect 296368 507134 296688 507218
rect 296368 506898 296410 507134
rect 296646 506898 296688 507134
rect 296368 506866 296688 506898
rect 327088 507454 327408 507486
rect 327088 507218 327130 507454
rect 327366 507218 327408 507454
rect 327088 507134 327408 507218
rect 327088 506898 327130 507134
rect 327366 506898 327408 507134
rect 327088 506866 327408 506898
rect 248459 501668 248525 501669
rect 248459 501604 248460 501668
rect 248524 501604 248525 501668
rect 248459 501603 248525 501604
rect 240114 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 240734 493774
rect 240114 493454 240734 493538
rect 240114 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 240734 493454
rect 240114 457774 240734 493218
rect 240114 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 240734 457774
rect 240114 457454 240734 457538
rect 240114 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 240734 457454
rect 240114 449580 240734 457218
rect 243834 497494 244454 501375
rect 243834 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 244454 497494
rect 243834 497174 244454 497258
rect 243834 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 244454 497174
rect 243834 461494 244454 496938
rect 243834 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 244454 461494
rect 243834 461174 244454 461258
rect 243834 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 244454 461174
rect 240288 439174 240608 439206
rect 240288 438938 240330 439174
rect 240566 438938 240608 439174
rect 240288 438854 240608 438938
rect 240288 438618 240330 438854
rect 240566 438618 240608 438854
rect 240288 438586 240608 438618
rect 236394 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 237014 418054
rect 236394 417734 237014 417818
rect 236394 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 237014 417734
rect 236394 382054 237014 417498
rect 243834 425494 244454 460938
rect 248462 452573 248522 501603
rect 253794 471454 254414 501375
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 248459 452572 248525 452573
rect 248459 452508 248460 452572
rect 248524 452508 248525 452572
rect 248459 452507 248525 452508
rect 243834 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 244454 425494
rect 243834 425174 244454 425258
rect 243834 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 244454 425174
rect 240288 403174 240608 403206
rect 240288 402938 240330 403174
rect 240566 402938 240608 403174
rect 240288 402854 240608 402938
rect 240288 402618 240330 402854
rect 240566 402618 240608 402854
rect 240288 402586 240608 402618
rect 236394 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 237014 382054
rect 236394 381734 237014 381818
rect 236394 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 237014 381734
rect 236394 346054 237014 381498
rect 243834 389494 244454 424938
rect 243834 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 244454 389494
rect 243834 389174 244454 389258
rect 243834 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 244454 389174
rect 240288 367174 240608 367206
rect 240288 366938 240330 367174
rect 240566 366938 240608 367174
rect 240288 366854 240608 366938
rect 240288 366618 240330 366854
rect 240566 366618 240608 366854
rect 240288 366586 240608 366618
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 236394 310054 237014 345498
rect 243834 353494 244454 388938
rect 243834 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 244454 353494
rect 243834 353174 244454 353258
rect 243834 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 244454 353174
rect 240288 331174 240608 331206
rect 240288 330938 240330 331174
rect 240566 330938 240608 331174
rect 240288 330854 240608 330938
rect 240288 330618 240330 330854
rect 240566 330618 240608 330854
rect 240288 330586 240608 330618
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 236394 274054 237014 309498
rect 243834 317494 244454 352938
rect 243834 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 244454 317494
rect 243834 317174 244454 317258
rect 243834 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 244454 317174
rect 240288 295174 240608 295206
rect 240288 294938 240330 295174
rect 240566 294938 240608 295174
rect 240288 294854 240608 294938
rect 240288 294618 240330 294854
rect 240566 294618 240608 294854
rect 240288 294586 240608 294618
rect 236394 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 237014 274054
rect 236394 273734 237014 273818
rect 236394 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 237014 273734
rect 236394 238054 237014 273498
rect 243834 281494 244454 316938
rect 243834 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 244454 281494
rect 243834 281174 244454 281258
rect 243834 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 244454 281174
rect 240288 259174 240608 259206
rect 240288 258938 240330 259174
rect 240566 258938 240608 259174
rect 240288 258854 240608 258938
rect 240288 258618 240330 258854
rect 240566 258618 240608 258854
rect 240288 258586 240608 258618
rect 236394 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 237014 238054
rect 236394 237734 237014 237818
rect 236394 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 237014 237734
rect 236394 202054 237014 237498
rect 236394 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 237014 202054
rect 236394 201734 237014 201818
rect 236394 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 237014 201734
rect 236394 166054 237014 201498
rect 236394 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 237014 166054
rect 236394 165734 237014 165818
rect 236394 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 237014 165734
rect 236394 130054 237014 165498
rect 236394 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 237014 130054
rect 236394 129734 237014 129818
rect 236394 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 237014 129734
rect 236394 105244 237014 129498
rect 240114 241774 240734 250068
rect 240114 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 240734 241774
rect 240114 241454 240734 241538
rect 240114 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 240734 241454
rect 240114 205774 240734 241218
rect 240114 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 240734 205774
rect 240114 205454 240734 205538
rect 240114 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 240734 205454
rect 240114 169774 240734 205218
rect 240114 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 240734 169774
rect 240114 169454 240734 169538
rect 240114 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 240734 169454
rect 240114 133774 240734 169218
rect 240114 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 240734 133774
rect 240114 133454 240734 133538
rect 240114 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 240734 133454
rect 240114 105244 240734 133218
rect 243834 245494 244454 280938
rect 243834 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 244454 245494
rect 243834 245174 244454 245258
rect 243834 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 244454 245174
rect 243834 209494 244454 244938
rect 243834 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 244454 209494
rect 243834 209174 244454 209258
rect 243834 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 244454 209174
rect 243834 173494 244454 208938
rect 243834 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 244454 173494
rect 243834 173174 244454 173258
rect 243834 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 244454 173174
rect 243834 137494 244454 172938
rect 243834 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 244454 137494
rect 243834 137174 244454 137258
rect 243834 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 244454 137174
rect 243834 105244 244454 136938
rect 253794 435454 254414 470898
rect 272394 490054 273014 501375
rect 272394 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 273014 490054
rect 272394 489734 273014 489818
rect 272394 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 273014 489734
rect 272394 454054 273014 489498
rect 272394 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 273014 454054
rect 272394 453734 273014 453818
rect 272394 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 273014 453734
rect 272394 451537 273014 453498
rect 276114 493774 276734 501375
rect 276114 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 276734 493774
rect 276114 493454 276734 493538
rect 276114 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 276734 493454
rect 276114 457774 276734 493218
rect 276114 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 276734 457774
rect 276114 457454 276734 457538
rect 276114 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 276734 457454
rect 276114 451537 276734 457218
rect 279834 497494 280454 501375
rect 279834 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 280454 497494
rect 279834 497174 280454 497258
rect 279834 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 280454 497174
rect 279834 461494 280454 496938
rect 279834 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 280454 461494
rect 279834 461174 280454 461258
rect 279834 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 280454 461174
rect 279834 451537 280454 460938
rect 308394 490054 309014 501375
rect 308394 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 309014 490054
rect 308394 489734 309014 489818
rect 308394 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 309014 489734
rect 308394 454054 309014 489498
rect 308394 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 309014 454054
rect 308394 453734 309014 453818
rect 308394 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 309014 453734
rect 308394 451537 309014 453498
rect 312114 493774 312734 501375
rect 312114 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 312734 493774
rect 312114 493454 312734 493538
rect 312114 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 312734 493454
rect 312114 457774 312734 493218
rect 312114 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 312734 457774
rect 312114 457454 312734 457538
rect 312114 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 312734 457454
rect 312114 451537 312734 457218
rect 315834 497494 316454 501375
rect 315834 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 316454 497494
rect 315834 497174 316454 497258
rect 315834 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 316454 497174
rect 315834 461494 316454 496938
rect 315834 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 316454 461494
rect 315834 461174 316454 461258
rect 315834 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 316454 461174
rect 315834 451537 316454 460938
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 451537 333854 478338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 451537 337574 482058
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 630334 341294 665778
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 342448 655174 342768 655206
rect 342448 654938 342490 655174
rect 342726 654938 342768 655174
rect 342448 654854 342768 654938
rect 342448 654618 342490 654854
rect 342726 654618 342768 654854
rect 342448 654586 342768 654618
rect 340674 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 341294 630334
rect 340674 630014 341294 630098
rect 340674 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 341294 630014
rect 340674 594334 341294 629778
rect 344394 634054 345014 669498
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 342448 619174 342768 619206
rect 342448 618938 342490 619174
rect 342726 618938 342768 619174
rect 342448 618854 342768 618938
rect 342448 618618 342490 618854
rect 342726 618618 342768 618854
rect 342448 618586 342768 618618
rect 340674 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 341294 594334
rect 340674 594014 341294 594098
rect 340674 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 341294 594014
rect 340674 558334 341294 593778
rect 344394 598054 345014 633498
rect 344394 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 345014 598054
rect 344394 597734 345014 597818
rect 344394 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 345014 597734
rect 342448 583174 342768 583206
rect 342448 582938 342490 583174
rect 342726 582938 342768 583174
rect 342448 582854 342768 582938
rect 342448 582618 342490 582854
rect 342726 582618 342768 582854
rect 342448 582586 342768 582618
rect 340674 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 341294 558334
rect 340674 558014 341294 558098
rect 340674 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 341294 558014
rect 340674 522334 341294 557778
rect 344394 562054 345014 597498
rect 344394 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 345014 562054
rect 344394 561734 345014 561818
rect 344394 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 345014 561734
rect 342448 547174 342768 547206
rect 342448 546938 342490 547174
rect 342726 546938 342768 547174
rect 342448 546854 342768 546938
rect 342448 546618 342490 546854
rect 342726 546618 342768 546854
rect 342448 546586 342768 546618
rect 340674 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 341294 522334
rect 340674 522014 341294 522098
rect 340674 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 341294 522014
rect 340674 486334 341294 521778
rect 344394 526054 345014 561498
rect 344394 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 345014 526054
rect 344394 525734 345014 525818
rect 344394 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 345014 525734
rect 342448 511174 342768 511206
rect 342448 510938 342490 511174
rect 342726 510938 342768 511174
rect 342448 510854 342768 510938
rect 342448 510618 342490 510854
rect 342726 510618 342768 510854
rect 342448 510586 342768 510618
rect 340674 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 341294 486334
rect 340674 486014 341294 486098
rect 340674 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 341294 486014
rect 340674 451537 341294 485778
rect 344394 490054 345014 525498
rect 344394 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 345014 490054
rect 344394 489734 345014 489818
rect 344394 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 345014 489734
rect 344394 454054 345014 489498
rect 344394 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 345014 454054
rect 344394 453734 345014 453818
rect 344394 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 345014 453734
rect 344394 451537 345014 453498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 348114 601774 348734 637218
rect 348114 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 348734 601774
rect 348114 601454 348734 601538
rect 348114 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 348734 601454
rect 348114 565774 348734 601218
rect 348114 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 348734 565774
rect 348114 565454 348734 565538
rect 348114 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 348734 565454
rect 348114 529774 348734 565218
rect 348114 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 348734 529774
rect 348114 529454 348734 529538
rect 348114 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 348734 529454
rect 348114 493774 348734 529218
rect 348114 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 348734 493774
rect 348114 493454 348734 493538
rect 348114 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 348734 493454
rect 348114 457774 348734 493218
rect 348114 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 348734 457774
rect 348114 457454 348734 457538
rect 348114 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 348734 457454
rect 348114 451537 348734 457218
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 357808 651454 358128 651486
rect 357808 651218 357850 651454
rect 358086 651218 358128 651454
rect 357808 651134 358128 651218
rect 357808 650898 357850 651134
rect 358086 650898 358128 651134
rect 357808 650866 358128 650898
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 605494 352454 640938
rect 357808 615454 358128 615486
rect 357808 615218 357850 615454
rect 358086 615218 358128 615454
rect 357808 615134 358128 615218
rect 357808 614898 357850 615134
rect 358086 614898 358128 615134
rect 357808 614866 358128 614898
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 351834 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 352454 605494
rect 351834 605174 352454 605258
rect 351834 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 352454 605174
rect 351834 569494 352454 604938
rect 357808 579454 358128 579486
rect 357808 579218 357850 579454
rect 358086 579218 358128 579454
rect 357808 579134 358128 579218
rect 357808 578898 357850 579134
rect 358086 578898 358128 579134
rect 357808 578866 358128 578898
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 351834 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 352454 569494
rect 351834 569174 352454 569258
rect 351834 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 352454 569174
rect 351834 533494 352454 568938
rect 357808 543454 358128 543486
rect 357808 543218 357850 543454
rect 358086 543218 358128 543454
rect 357808 543134 358128 543218
rect 357808 542898 357850 543134
rect 358086 542898 358128 543134
rect 357808 542866 358128 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 351834 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 352454 533494
rect 351834 533174 352454 533258
rect 351834 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 352454 533174
rect 351834 497494 352454 532938
rect 357808 507454 358128 507486
rect 357808 507218 357850 507454
rect 358086 507218 358128 507454
rect 357808 507134 358128 507218
rect 357808 506898 357850 507134
rect 358086 506898 358128 507134
rect 357808 506866 358128 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 351834 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 352454 497494
rect 351834 497174 352454 497258
rect 351834 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 352454 497174
rect 351834 461494 352454 496938
rect 351834 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 352454 461494
rect 351834 461174 352454 461258
rect 351834 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 352454 461174
rect 351834 451537 352454 460938
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 451537 362414 470898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 451537 366134 474618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372659 682140 372725 682141
rect 372659 682076 372660 682140
rect 372724 682076 372725 682140
rect 372659 682075 372725 682076
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 372662 494869 372722 682075
rect 372954 679452 373574 698058
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 374131 682684 374197 682685
rect 374131 682620 374132 682684
rect 374196 682620 374197 682684
rect 374131 682619 374197 682620
rect 373763 682276 373829 682277
rect 373763 682212 373764 682276
rect 373828 682212 373829 682276
rect 373763 682211 373829 682212
rect 373168 655174 373488 655206
rect 373168 654938 373210 655174
rect 373446 654938 373488 655174
rect 373168 654854 373488 654938
rect 373168 654618 373210 654854
rect 373446 654618 373488 654854
rect 373168 654586 373488 654618
rect 373168 619174 373488 619206
rect 373168 618938 373210 619174
rect 373446 618938 373488 619174
rect 373168 618854 373488 618938
rect 373168 618618 373210 618854
rect 373446 618618 373488 618854
rect 373168 618586 373488 618618
rect 373168 583174 373488 583206
rect 373168 582938 373210 583174
rect 373446 582938 373488 583174
rect 373168 582854 373488 582938
rect 373168 582618 373210 582854
rect 373446 582618 373488 582854
rect 373168 582586 373488 582618
rect 373168 547174 373488 547206
rect 373168 546938 373210 547174
rect 373446 546938 373488 547174
rect 373168 546854 373488 546938
rect 373168 546618 373210 546854
rect 373446 546618 373488 546854
rect 373168 546586 373488 546618
rect 373168 511174 373488 511206
rect 373168 510938 373210 511174
rect 373446 510938 373488 511174
rect 373168 510854 373488 510938
rect 373168 510618 373210 510854
rect 373446 510618 373488 510854
rect 373168 510586 373488 510618
rect 372659 494868 372725 494869
rect 372659 494804 372660 494868
rect 372724 494804 372725 494868
rect 372659 494803 372725 494804
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 271008 439174 271328 439206
rect 271008 438938 271050 439174
rect 271286 438938 271328 439174
rect 271008 438854 271328 438938
rect 271008 438618 271050 438854
rect 271286 438618 271328 438854
rect 271008 438586 271328 438618
rect 301728 439174 302048 439206
rect 301728 438938 301770 439174
rect 302006 438938 302048 439174
rect 301728 438854 302048 438938
rect 301728 438618 301770 438854
rect 302006 438618 302048 438854
rect 301728 438586 302048 438618
rect 332448 439174 332768 439206
rect 332448 438938 332490 439174
rect 332726 438938 332768 439174
rect 332448 438854 332768 438938
rect 332448 438618 332490 438854
rect 332726 438618 332768 438854
rect 332448 438586 332768 438618
rect 363168 439174 363488 439206
rect 363168 438938 363210 439174
rect 363446 438938 363488 439174
rect 363168 438854 363488 438938
rect 363168 438618 363210 438854
rect 363446 438618 363488 438854
rect 363168 438586 363488 438618
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 255648 435454 255968 435486
rect 255648 435218 255690 435454
rect 255926 435218 255968 435454
rect 255648 435134 255968 435218
rect 255648 434898 255690 435134
rect 255926 434898 255968 435134
rect 255648 434866 255968 434898
rect 286368 435454 286688 435486
rect 286368 435218 286410 435454
rect 286646 435218 286688 435454
rect 286368 435134 286688 435218
rect 286368 434898 286410 435134
rect 286646 434898 286688 435134
rect 286368 434866 286688 434898
rect 317088 435454 317408 435486
rect 317088 435218 317130 435454
rect 317366 435218 317408 435454
rect 317088 435134 317408 435218
rect 317088 434898 317130 435134
rect 317366 434898 317408 435134
rect 317088 434866 317408 434898
rect 347808 435454 348128 435486
rect 347808 435218 347850 435454
rect 348086 435218 348128 435454
rect 347808 435134 348128 435218
rect 347808 434898 347850 435134
rect 348086 434898 348128 435134
rect 347808 434866 348128 434898
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 271008 403174 271328 403206
rect 271008 402938 271050 403174
rect 271286 402938 271328 403174
rect 271008 402854 271328 402938
rect 271008 402618 271050 402854
rect 271286 402618 271328 402854
rect 271008 402586 271328 402618
rect 301728 403174 302048 403206
rect 301728 402938 301770 403174
rect 302006 402938 302048 403174
rect 301728 402854 302048 402938
rect 301728 402618 301770 402854
rect 302006 402618 302048 402854
rect 301728 402586 302048 402618
rect 332448 403174 332768 403206
rect 332448 402938 332490 403174
rect 332726 402938 332768 403174
rect 332448 402854 332768 402938
rect 332448 402618 332490 402854
rect 332726 402618 332768 402854
rect 332448 402586 332768 402618
rect 363168 403174 363488 403206
rect 363168 402938 363210 403174
rect 363446 402938 363488 403174
rect 363168 402854 363488 402938
rect 363168 402618 363210 402854
rect 363446 402618 363488 402854
rect 363168 402586 363488 402618
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 255648 399454 255968 399486
rect 255648 399218 255690 399454
rect 255926 399218 255968 399454
rect 255648 399134 255968 399218
rect 255648 398898 255690 399134
rect 255926 398898 255968 399134
rect 255648 398866 255968 398898
rect 286368 399454 286688 399486
rect 286368 399218 286410 399454
rect 286646 399218 286688 399454
rect 286368 399134 286688 399218
rect 286368 398898 286410 399134
rect 286646 398898 286688 399134
rect 286368 398866 286688 398898
rect 317088 399454 317408 399486
rect 317088 399218 317130 399454
rect 317366 399218 317408 399454
rect 317088 399134 317408 399218
rect 317088 398898 317130 399134
rect 317366 398898 317408 399134
rect 317088 398866 317408 398898
rect 347808 399454 348128 399486
rect 347808 399218 347850 399454
rect 348086 399218 348128 399454
rect 347808 399134 348128 399218
rect 347808 398898 347850 399134
rect 348086 398898 348128 399134
rect 347808 398866 348128 398898
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 271008 367174 271328 367206
rect 271008 366938 271050 367174
rect 271286 366938 271328 367174
rect 271008 366854 271328 366938
rect 271008 366618 271050 366854
rect 271286 366618 271328 366854
rect 271008 366586 271328 366618
rect 301728 367174 302048 367206
rect 301728 366938 301770 367174
rect 302006 366938 302048 367174
rect 301728 366854 302048 366938
rect 301728 366618 301770 366854
rect 302006 366618 302048 366854
rect 301728 366586 302048 366618
rect 332448 367174 332768 367206
rect 332448 366938 332490 367174
rect 332726 366938 332768 367174
rect 332448 366854 332768 366938
rect 332448 366618 332490 366854
rect 332726 366618 332768 366854
rect 332448 366586 332768 366618
rect 363168 367174 363488 367206
rect 363168 366938 363210 367174
rect 363446 366938 363488 367174
rect 363168 366854 363488 366938
rect 363168 366618 363210 366854
rect 363446 366618 363488 366854
rect 363168 366586 363488 366618
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 255648 363454 255968 363486
rect 255648 363218 255690 363454
rect 255926 363218 255968 363454
rect 255648 363134 255968 363218
rect 255648 362898 255690 363134
rect 255926 362898 255968 363134
rect 255648 362866 255968 362898
rect 286368 363454 286688 363486
rect 286368 363218 286410 363454
rect 286646 363218 286688 363454
rect 286368 363134 286688 363218
rect 286368 362898 286410 363134
rect 286646 362898 286688 363134
rect 286368 362866 286688 362898
rect 317088 363454 317408 363486
rect 317088 363218 317130 363454
rect 317366 363218 317408 363454
rect 317088 363134 317408 363218
rect 317088 362898 317130 363134
rect 317366 362898 317408 363134
rect 317088 362866 317408 362898
rect 347808 363454 348128 363486
rect 347808 363218 347850 363454
rect 348086 363218 348128 363454
rect 347808 363134 348128 363218
rect 347808 362898 347850 363134
rect 348086 362898 348128 363134
rect 347808 362866 348128 362898
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 271008 331174 271328 331206
rect 271008 330938 271050 331174
rect 271286 330938 271328 331174
rect 271008 330854 271328 330938
rect 271008 330618 271050 330854
rect 271286 330618 271328 330854
rect 271008 330586 271328 330618
rect 301728 331174 302048 331206
rect 301728 330938 301770 331174
rect 302006 330938 302048 331174
rect 301728 330854 302048 330938
rect 301728 330618 301770 330854
rect 302006 330618 302048 330854
rect 301728 330586 302048 330618
rect 332448 331174 332768 331206
rect 332448 330938 332490 331174
rect 332726 330938 332768 331174
rect 332448 330854 332768 330938
rect 332448 330618 332490 330854
rect 332726 330618 332768 330854
rect 332448 330586 332768 330618
rect 363168 331174 363488 331206
rect 363168 330938 363210 331174
rect 363446 330938 363488 331174
rect 363168 330854 363488 330938
rect 363168 330618 363210 330854
rect 363446 330618 363488 330854
rect 363168 330586 363488 330618
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 255648 327454 255968 327486
rect 255648 327218 255690 327454
rect 255926 327218 255968 327454
rect 255648 327134 255968 327218
rect 255648 326898 255690 327134
rect 255926 326898 255968 327134
rect 255648 326866 255968 326898
rect 286368 327454 286688 327486
rect 286368 327218 286410 327454
rect 286646 327218 286688 327454
rect 286368 327134 286688 327218
rect 286368 326898 286410 327134
rect 286646 326898 286688 327134
rect 286368 326866 286688 326898
rect 317088 327454 317408 327486
rect 317088 327218 317130 327454
rect 317366 327218 317408 327454
rect 317088 327134 317408 327218
rect 317088 326898 317130 327134
rect 317366 326898 317408 327134
rect 317088 326866 317408 326898
rect 347808 327454 348128 327486
rect 347808 327218 347850 327454
rect 348086 327218 348128 327454
rect 347808 327134 348128 327218
rect 347808 326898 347850 327134
rect 348086 326898 348128 327134
rect 347808 326866 348128 326898
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 271008 295174 271328 295206
rect 271008 294938 271050 295174
rect 271286 294938 271328 295174
rect 271008 294854 271328 294938
rect 271008 294618 271050 294854
rect 271286 294618 271328 294854
rect 271008 294586 271328 294618
rect 301728 295174 302048 295206
rect 301728 294938 301770 295174
rect 302006 294938 302048 295174
rect 301728 294854 302048 294938
rect 301728 294618 301770 294854
rect 302006 294618 302048 294854
rect 301728 294586 302048 294618
rect 332448 295174 332768 295206
rect 332448 294938 332490 295174
rect 332726 294938 332768 295174
rect 332448 294854 332768 294938
rect 332448 294618 332490 294854
rect 332726 294618 332768 294854
rect 332448 294586 332768 294618
rect 363168 295174 363488 295206
rect 363168 294938 363210 295174
rect 363446 294938 363488 295174
rect 363168 294854 363488 294938
rect 363168 294618 363210 294854
rect 363446 294618 363488 294854
rect 363168 294586 363488 294618
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 255648 291454 255968 291486
rect 255648 291218 255690 291454
rect 255926 291218 255968 291454
rect 255648 291134 255968 291218
rect 255648 290898 255690 291134
rect 255926 290898 255968 291134
rect 255648 290866 255968 290898
rect 286368 291454 286688 291486
rect 286368 291218 286410 291454
rect 286646 291218 286688 291454
rect 286368 291134 286688 291218
rect 286368 290898 286410 291134
rect 286646 290898 286688 291134
rect 286368 290866 286688 290898
rect 317088 291454 317408 291486
rect 317088 291218 317130 291454
rect 317366 291218 317408 291454
rect 317088 291134 317408 291218
rect 317088 290898 317130 291134
rect 317366 290898 317408 291134
rect 317088 290866 317408 290898
rect 347808 291454 348128 291486
rect 347808 291218 347850 291454
rect 348086 291218 348128 291454
rect 347808 291134 348128 291218
rect 347808 290898 347850 291134
rect 348086 290898 348128 291134
rect 347808 290866 348128 290898
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 271008 259174 271328 259206
rect 271008 258938 271050 259174
rect 271286 258938 271328 259174
rect 271008 258854 271328 258938
rect 271008 258618 271050 258854
rect 271286 258618 271328 258854
rect 271008 258586 271328 258618
rect 301728 259174 302048 259206
rect 301728 258938 301770 259174
rect 302006 258938 302048 259174
rect 301728 258854 302048 258938
rect 301728 258618 301770 258854
rect 302006 258618 302048 258854
rect 301728 258586 302048 258618
rect 332448 259174 332768 259206
rect 332448 258938 332490 259174
rect 332726 258938 332768 259174
rect 332448 258854 332768 258938
rect 332448 258618 332490 258854
rect 332726 258618 332768 258854
rect 332448 258586 332768 258618
rect 363168 259174 363488 259206
rect 363168 258938 363210 259174
rect 363446 258938 363488 259174
rect 363168 258854 363488 258938
rect 363168 258618 363210 258854
rect 363446 258618 363488 258854
rect 363168 258586 363488 258618
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 255648 255454 255968 255486
rect 255648 255218 255690 255454
rect 255926 255218 255968 255454
rect 255648 255134 255968 255218
rect 255648 254898 255690 255134
rect 255926 254898 255968 255134
rect 255648 254866 255968 254898
rect 286368 255454 286688 255486
rect 286368 255218 286410 255454
rect 286646 255218 286688 255454
rect 286368 255134 286688 255218
rect 286368 254898 286410 255134
rect 286646 254898 286688 255134
rect 286368 254866 286688 254898
rect 317088 255454 317408 255486
rect 317088 255218 317130 255454
rect 317366 255218 317408 255454
rect 317088 255134 317408 255218
rect 317088 254898 317130 255134
rect 317366 254898 317408 255134
rect 317088 254866 317408 254898
rect 347808 255454 348128 255486
rect 347808 255218 347850 255454
rect 348086 255218 348128 255454
rect 347808 255134 348128 255218
rect 347808 254898 347850 255134
rect 348086 254898 348128 255134
rect 347808 254866 348128 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 105244 254414 110898
rect 257514 223174 258134 249743
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 105244 258134 114618
rect 261234 226894 261854 249743
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 105244 261854 118338
rect 264954 230614 265574 249743
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 105244 265574 122058
rect 268674 234334 269294 249743
rect 268674 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 269294 234334
rect 268674 234014 269294 234098
rect 268674 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 269294 234014
rect 268674 198334 269294 233778
rect 268674 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 269294 198334
rect 268674 198014 269294 198098
rect 268674 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 269294 198014
rect 268674 162334 269294 197778
rect 268674 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 269294 162334
rect 268674 162014 269294 162098
rect 268674 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 269294 162014
rect 268674 126334 269294 161778
rect 268674 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 269294 126334
rect 268674 126014 269294 126098
rect 268674 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 269294 126014
rect 268674 105244 269294 125778
rect 272394 238054 273014 249743
rect 272394 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 273014 238054
rect 272394 237734 273014 237818
rect 272394 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 273014 237734
rect 272394 202054 273014 237498
rect 272394 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 273014 202054
rect 272394 201734 273014 201818
rect 272394 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 273014 201734
rect 272394 166054 273014 201498
rect 272394 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 273014 166054
rect 272394 165734 273014 165818
rect 272394 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 273014 165734
rect 272394 130054 273014 165498
rect 272394 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 273014 130054
rect 272394 129734 273014 129818
rect 272394 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 273014 129734
rect 272394 105244 273014 129498
rect 276114 241774 276734 249743
rect 276114 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 276734 241774
rect 276114 241454 276734 241538
rect 276114 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 276734 241454
rect 276114 205774 276734 241218
rect 276114 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 276734 205774
rect 276114 205454 276734 205538
rect 276114 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 276734 205454
rect 276114 169774 276734 205218
rect 276114 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 276734 169774
rect 276114 169454 276734 169538
rect 276114 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 276734 169454
rect 276114 133774 276734 169218
rect 276114 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 276734 133774
rect 276114 133454 276734 133538
rect 276114 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 276734 133454
rect 276114 105244 276734 133218
rect 279834 245494 280454 249743
rect 279834 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 280454 245494
rect 279834 245174 280454 245258
rect 279834 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 280454 245174
rect 279834 209494 280454 244938
rect 279834 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 280454 209494
rect 279834 209174 280454 209258
rect 279834 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 280454 209174
rect 279834 173494 280454 208938
rect 279834 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 280454 173494
rect 279834 173174 280454 173258
rect 279834 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 280454 173174
rect 279834 137494 280454 172938
rect 279834 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 280454 137494
rect 279834 137174 280454 137258
rect 279834 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 280454 137174
rect 279834 105244 280454 136938
rect 289794 219454 290414 249743
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 105244 290414 110898
rect 293514 223174 294134 249743
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 105244 294134 114618
rect 297234 226894 297854 249743
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 105244 297854 118338
rect 300954 230614 301574 249743
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 105244 301574 122058
rect 304674 234334 305294 249743
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 304674 198334 305294 233778
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 304674 162334 305294 197778
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 304674 126334 305294 161778
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 304674 105244 305294 125778
rect 308394 238054 309014 249743
rect 308394 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 309014 238054
rect 308394 237734 309014 237818
rect 308394 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 309014 237734
rect 308394 202054 309014 237498
rect 308394 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 309014 202054
rect 308394 201734 309014 201818
rect 308394 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 309014 201734
rect 308394 166054 309014 201498
rect 308394 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 309014 166054
rect 308394 165734 309014 165818
rect 308394 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 309014 165734
rect 308394 130054 309014 165498
rect 308394 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 309014 130054
rect 308394 129734 309014 129818
rect 308394 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 309014 129734
rect 308394 105244 309014 129498
rect 312114 241774 312734 249743
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 312114 205774 312734 241218
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 312114 169774 312734 205218
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 312114 133774 312734 169218
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 312114 105244 312734 133218
rect 315834 245494 316454 249743
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 315834 209494 316454 244938
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 315834 173494 316454 208938
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 315834 105244 316454 136938
rect 325794 219454 326414 249743
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 105244 326414 110898
rect 329514 223174 330134 249743
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 105244 330134 114618
rect 333234 226894 333854 249743
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 105244 333854 118338
rect 336954 230614 337574 249743
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 105244 337574 122058
rect 340674 234334 341294 249743
rect 340674 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 341294 234334
rect 340674 234014 341294 234098
rect 340674 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 341294 234014
rect 340674 198334 341294 233778
rect 340674 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 341294 198334
rect 340674 198014 341294 198098
rect 340674 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 341294 198014
rect 340674 162334 341294 197778
rect 340674 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 341294 162334
rect 340674 162014 341294 162098
rect 340674 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 341294 162014
rect 340674 126334 341294 161778
rect 340674 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 341294 126334
rect 340674 126014 341294 126098
rect 340674 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 341294 126014
rect 340674 105244 341294 125778
rect 344394 238054 345014 249743
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 344394 202054 345014 237498
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 344394 166054 345014 201498
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 344394 130054 345014 165498
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 344394 105244 345014 129498
rect 348114 241774 348734 249743
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 348114 169774 348734 205218
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 348114 133774 348734 169218
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 348114 105244 348734 133218
rect 351834 245494 352454 249743
rect 357203 247212 357269 247213
rect 357203 247148 357204 247212
rect 357268 247148 357269 247212
rect 357203 247147 357269 247148
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 351834 173494 352454 208938
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 350947 106180 351013 106181
rect 350947 106116 350948 106180
rect 351012 106116 351013 106180
rect 350947 106115 351013 106116
rect 350950 103530 351010 106115
rect 351834 105244 352454 136938
rect 350840 103470 351010 103530
rect 350840 103202 350900 103470
rect 207834 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 208454 101494
rect 207834 101174 208454 101258
rect 207834 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 208454 101174
rect 207834 65494 208454 100938
rect 220272 79174 220620 79206
rect 220272 78938 220328 79174
rect 220564 78938 220620 79174
rect 220272 78854 220620 78938
rect 220272 78618 220328 78854
rect 220564 78618 220620 78854
rect 220272 78586 220620 78618
rect 356000 79174 356348 79206
rect 356000 78938 356056 79174
rect 356292 78938 356348 79174
rect 356000 78854 356348 78938
rect 356000 78618 356056 78854
rect 356292 78618 356348 78854
rect 356000 78586 356348 78618
rect 220952 75454 221300 75486
rect 220952 75218 221008 75454
rect 221244 75218 221300 75454
rect 220952 75134 221300 75218
rect 220952 74898 221008 75134
rect 221244 74898 221300 75134
rect 220952 74866 221300 74898
rect 355320 75454 355668 75486
rect 355320 75218 355376 75454
rect 355612 75218 355668 75454
rect 355320 75134 355668 75218
rect 355320 74898 355376 75134
rect 355612 74898 355668 75134
rect 355320 74866 355668 74898
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 207834 29494 208454 64938
rect 220272 43174 220620 43206
rect 220272 42938 220328 43174
rect 220564 42938 220620 43174
rect 220272 42854 220620 42938
rect 220272 42618 220328 42854
rect 220564 42618 220620 42854
rect 220272 42586 220620 42618
rect 356000 43174 356348 43206
rect 356000 42938 356056 43174
rect 356292 42938 356348 43174
rect 356000 42854 356348 42938
rect 356000 42618 356056 42854
rect 356292 42618 356348 42854
rect 356000 42586 356348 42618
rect 220952 39454 221300 39486
rect 220952 39218 221008 39454
rect 221244 39218 221300 39454
rect 220952 39134 221300 39218
rect 220952 38898 221008 39134
rect 221244 38898 221300 39134
rect 220952 38866 221300 38898
rect 355320 39454 355668 39486
rect 355320 39218 355376 39454
rect 355612 39218 355668 39454
rect 355320 39134 355668 39218
rect 355320 38898 355376 39134
rect 355612 38898 355668 39134
rect 355320 38866 355668 38898
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 236056 19410 236116 20060
rect 237144 19410 237204 20060
rect 238232 19410 238292 20060
rect 239592 19682 239652 20060
rect 240544 19682 240604 20060
rect 241768 19682 241828 20060
rect 243128 19682 243188 20060
rect 239592 19622 239690 19682
rect 240544 19622 240610 19682
rect 235950 19350 236116 19410
rect 237054 19350 237204 19410
rect 238158 19350 238292 19410
rect 235950 18597 236010 19350
rect 237054 18733 237114 19350
rect 238158 18869 238218 19350
rect 239630 19141 239690 19622
rect 240550 19277 240610 19622
rect 241654 19622 241828 19682
rect 243126 19622 243188 19682
rect 244216 19682 244276 20060
rect 245440 19682 245500 20060
rect 246528 19682 246588 20060
rect 247616 19682 247676 20060
rect 248296 19682 248356 20060
rect 248704 19682 248764 20060
rect 244216 19622 244290 19682
rect 240547 19276 240613 19277
rect 240547 19212 240548 19276
rect 240612 19212 240613 19276
rect 240547 19211 240613 19212
rect 239627 19140 239693 19141
rect 239627 19076 239628 19140
rect 239692 19076 239693 19140
rect 239627 19075 239693 19076
rect 241654 19005 241714 19622
rect 241651 19004 241717 19005
rect 241651 18940 241652 19004
rect 241716 18940 241717 19004
rect 241651 18939 241717 18940
rect 238155 18868 238221 18869
rect 238155 18804 238156 18868
rect 238220 18804 238221 18868
rect 238155 18803 238221 18804
rect 237051 18732 237117 18733
rect 237051 18668 237052 18732
rect 237116 18668 237117 18732
rect 237051 18667 237117 18668
rect 243126 18597 243186 19622
rect 244230 19277 244290 19622
rect 245334 19622 245500 19682
rect 246438 19622 246588 19682
rect 247542 19622 247676 19682
rect 248278 19622 248356 19682
rect 248646 19622 248764 19682
rect 250064 19682 250124 20060
rect 250744 19682 250804 20060
rect 251288 19682 251348 20060
rect 252376 19682 252436 20060
rect 253464 19682 253524 20060
rect 250064 19622 250178 19682
rect 245334 19277 245394 19622
rect 246438 19277 246498 19622
rect 244227 19276 244293 19277
rect 244227 19212 244228 19276
rect 244292 19212 244293 19276
rect 244227 19211 244293 19212
rect 245331 19276 245397 19277
rect 245331 19212 245332 19276
rect 245396 19212 245397 19276
rect 245331 19211 245397 19212
rect 246435 19276 246501 19277
rect 246435 19212 246436 19276
rect 246500 19212 246501 19276
rect 246435 19211 246501 19212
rect 247542 19005 247602 19622
rect 248278 19141 248338 19622
rect 248275 19140 248341 19141
rect 248275 19076 248276 19140
rect 248340 19076 248341 19140
rect 248275 19075 248341 19076
rect 247539 19004 247605 19005
rect 247539 18940 247540 19004
rect 247604 18940 247605 19004
rect 247539 18939 247605 18940
rect 235947 18596 236013 18597
rect 235947 18532 235948 18596
rect 236012 18532 236013 18596
rect 235947 18531 236013 18532
rect 243123 18596 243189 18597
rect 243123 18532 243124 18596
rect 243188 18532 243189 18596
rect 243123 18531 243189 18532
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 3454 218414 18064
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 7174 222134 18064
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 10894 225854 18064
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 14614 229574 18064
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18023 233294 18064
rect 232674 17787 232706 18023
rect 232942 17787 233026 18023
rect 233262 17787 233294 18023
rect 232674 -4186 233294 17787
rect 248646 17373 248706 19622
rect 250118 19141 250178 19622
rect 250670 19622 250804 19682
rect 251222 19622 251348 19682
rect 252326 19622 252436 19682
rect 253430 19622 253524 19682
rect 253600 19682 253660 20060
rect 254552 19682 254612 20060
rect 255912 19682 255972 20060
rect 253600 19622 253674 19682
rect 250115 19140 250181 19141
rect 250115 19076 250116 19140
rect 250180 19076 250181 19140
rect 250115 19075 250181 19076
rect 250670 19005 250730 19622
rect 250667 19004 250733 19005
rect 250667 18940 250668 19004
rect 250732 18940 250733 19004
rect 250667 18939 250733 18940
rect 248643 17372 248709 17373
rect 248643 17308 248644 17372
rect 248708 17308 248709 17372
rect 248643 17307 248709 17308
rect 251222 17101 251282 19622
rect 252326 18869 252386 19622
rect 252323 18868 252389 18869
rect 252323 18804 252324 18868
rect 252388 18804 252389 18868
rect 252323 18803 252389 18804
rect 253430 17509 253490 19622
rect 253614 18869 253674 19622
rect 254534 19622 254612 19682
rect 255822 19622 255972 19682
rect 253611 18868 253677 18869
rect 253611 18804 253612 18868
rect 253676 18804 253677 18868
rect 253611 18803 253677 18804
rect 253427 17508 253493 17509
rect 253427 17444 253428 17508
rect 253492 17444 253493 17508
rect 253427 17443 253493 17444
rect 251219 17100 251285 17101
rect 251219 17036 251220 17100
rect 251284 17036 251285 17100
rect 251219 17035 251285 17036
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 253794 3454 254414 18064
rect 254534 17645 254594 19622
rect 254531 17644 254597 17645
rect 254531 17580 254532 17644
rect 254596 17580 254597 17644
rect 254531 17579 254597 17580
rect 255822 17373 255882 19622
rect 256048 19410 256108 20060
rect 257000 19682 257060 20060
rect 256006 19350 256108 19410
rect 256926 19622 257060 19682
rect 256006 18733 256066 19350
rect 256003 18732 256069 18733
rect 256003 18668 256004 18732
rect 256068 18668 256069 18732
rect 256003 18667 256069 18668
rect 256926 17373 256986 19622
rect 258088 19410 258148 20060
rect 258496 19410 258556 20060
rect 258088 19350 258274 19410
rect 255819 17372 255885 17373
rect 255819 17308 255820 17372
rect 255884 17308 255885 17372
rect 255819 17307 255885 17308
rect 256923 17372 256989 17373
rect 256923 17308 256924 17372
rect 256988 17308 256989 17372
rect 256923 17307 256989 17308
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 7174 258134 17940
rect 258214 17370 258274 19350
rect 258398 19350 258556 19410
rect 259448 19410 259508 20060
rect 260672 19410 260732 20060
rect 261080 19410 261140 20060
rect 259448 19350 259562 19410
rect 258398 18733 258458 19350
rect 258395 18732 258461 18733
rect 258395 18668 258396 18732
rect 258460 18668 258461 18732
rect 258395 18667 258461 18668
rect 259502 17509 259562 19350
rect 260606 19350 260732 19410
rect 260974 19350 261140 19410
rect 263528 19410 263588 20060
rect 265976 19410 266036 20060
rect 263528 19350 263610 19410
rect 260606 17645 260666 19350
rect 260974 17645 261034 19350
rect 260603 17644 260669 17645
rect 260603 17580 260604 17644
rect 260668 17580 260669 17644
rect 260603 17579 260669 17580
rect 260971 17644 261037 17645
rect 260971 17580 260972 17644
rect 261036 17580 261037 17644
rect 260971 17579 261037 17580
rect 259499 17508 259565 17509
rect 259499 17444 259500 17508
rect 259564 17444 259565 17508
rect 259499 17443 259565 17444
rect 258395 17372 258461 17373
rect 258395 17370 258396 17372
rect 258214 17310 258396 17370
rect 258395 17308 258396 17310
rect 258460 17308 258461 17372
rect 258395 17307 258461 17308
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 10894 261854 17940
rect 263550 17781 263610 19350
rect 265942 19350 266036 19410
rect 268288 19410 268348 20060
rect 271008 19410 271068 20060
rect 273592 19410 273652 20060
rect 268288 19350 268394 19410
rect 263547 17780 263613 17781
rect 263547 17716 263548 17780
rect 263612 17716 263613 17780
rect 263547 17715 263613 17716
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 17940
rect 265942 17781 266002 19350
rect 268334 17917 268394 19350
rect 270910 19350 271068 19410
rect 273486 19350 273652 19410
rect 276040 19410 276100 20060
rect 278488 19410 278548 20060
rect 280936 19410 280996 20060
rect 283520 19410 283580 20060
rect 285968 19549 286028 20060
rect 285965 19548 286031 19549
rect 285965 19484 285966 19548
rect 286030 19484 286031 19548
rect 285965 19483 286031 19484
rect 276040 19350 276122 19410
rect 268331 17916 268397 17917
rect 268331 17852 268332 17916
rect 268396 17852 268397 17916
rect 268331 17851 268397 17852
rect 265939 17780 266005 17781
rect 265939 17716 265940 17780
rect 266004 17716 266005 17780
rect 265939 17715 266005 17716
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 -4186 269294 17940
rect 270910 17645 270970 19350
rect 273486 17917 273546 19350
rect 273483 17916 273549 17917
rect 273483 17852 273484 17916
rect 273548 17852 273549 17916
rect 273483 17851 273549 17852
rect 270907 17644 270973 17645
rect 270907 17580 270908 17644
rect 270972 17580 270973 17644
rect 270907 17579 270973 17580
rect 276062 17237 276122 19350
rect 277166 19350 278548 19410
rect 280846 19350 280996 19410
rect 283422 19350 283580 19410
rect 277166 17917 277226 19350
rect 280846 17917 280906 19350
rect 277163 17916 277229 17917
rect 277163 17852 277164 17916
rect 277228 17852 277229 17916
rect 277163 17851 277229 17852
rect 280843 17916 280909 17917
rect 280843 17852 280844 17916
rect 280908 17852 280909 17916
rect 280843 17851 280909 17852
rect 283422 17237 283482 19350
rect 276059 17236 276125 17237
rect 276059 17172 276060 17236
rect 276124 17172 276125 17236
rect 276059 17171 276125 17172
rect 283419 17236 283485 17237
rect 283419 17172 283420 17236
rect 283484 17172 283485 17236
rect 283419 17171 283485 17172
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 289794 3454 290414 18064
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 7174 294134 17940
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 10894 297854 18064
rect 304674 18023 305294 18064
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 17940
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 17787 304706 18023
rect 304942 17787 305026 18023
rect 305262 17787 305294 18023
rect 304674 -4186 305294 17787
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 325794 3454 326414 17940
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 7174 330134 18064
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 10894 333854 18064
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 14614 337574 18064
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 18023 341294 18064
rect 340674 17787 340706 18023
rect 340942 17787 341026 18023
rect 341262 17787 341294 18023
rect 340674 -4186 341294 17787
rect 357206 7717 357266 247147
rect 359963 247076 360029 247077
rect 359963 247012 359964 247076
rect 360028 247012 360029 247076
rect 359963 247011 360029 247012
rect 357203 7716 357269 7717
rect 357203 7652 357204 7716
rect 357268 7652 357269 7716
rect 357203 7651 357269 7652
rect 359966 7581 360026 247011
rect 361794 219454 362414 249743
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 359963 7580 360029 7581
rect 359963 7516 359964 7580
rect 360028 7516 360029 7580
rect 359963 7515 360029 7516
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 223174 366134 249743
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 482614 373574 500068
rect 373766 494733 373826 682211
rect 374134 495005 374194 682619
rect 375419 682548 375485 682549
rect 375419 682484 375420 682548
rect 375484 682484 375485 682548
rect 375419 682483 375485 682484
rect 374499 584356 374565 584357
rect 374499 584292 374500 584356
rect 374564 584292 374565 584356
rect 374499 584291 374565 584292
rect 374131 495004 374197 495005
rect 374131 494940 374132 495004
rect 374196 494940 374197 495004
rect 374131 494939 374197 494940
rect 373763 494732 373829 494733
rect 373763 494668 373764 494732
rect 373828 494668 373829 494732
rect 373763 494667 373829 494668
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 374502 452573 374562 584291
rect 375422 500717 375482 682483
rect 376674 666334 377294 708122
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 378179 682412 378245 682413
rect 378179 682348 378180 682412
rect 378244 682348 378245 682412
rect 378179 682347 378245 682348
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376339 585716 376405 585717
rect 376339 585652 376340 585716
rect 376404 585652 376405 585716
rect 376339 585651 376405 585652
rect 375419 500716 375485 500717
rect 375419 500652 375420 500716
rect 375484 500652 375485 500716
rect 375419 500651 375485 500652
rect 376342 452573 376402 585651
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 378182 497589 378242 682347
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 378179 497588 378245 497589
rect 378179 497524 378180 497588
rect 378244 497524 378245 497588
rect 378179 497523 378245 497524
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 374499 452572 374565 452573
rect 374499 452508 374500 452572
rect 374564 452508 374565 452572
rect 374499 452507 374565 452508
rect 376339 452572 376405 452573
rect 376339 452508 376340 452572
rect 376404 452508 376405 452572
rect 376339 452507 376405 452508
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 378528 435454 378848 435486
rect 378528 435218 378570 435454
rect 378806 435218 378848 435454
rect 378528 435134 378848 435218
rect 378528 434898 378570 435134
rect 378806 434898 378848 435134
rect 378528 434866 378848 434898
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 378528 399454 378848 399486
rect 378528 399218 378570 399454
rect 378806 399218 378848 399454
rect 378528 399134 378848 399218
rect 378528 398898 378570 399134
rect 378806 398898 378848 399134
rect 378528 398866 378848 398898
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 378528 363454 378848 363486
rect 378528 363218 378570 363454
rect 378806 363218 378848 363454
rect 378528 363134 378848 363218
rect 378528 362898 378570 363134
rect 378806 362898 378848 363134
rect 378528 362866 378848 362898
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 378528 327454 378848 327486
rect 378528 327218 378570 327454
rect 378806 327218 378848 327454
rect 378528 327134 378848 327218
rect 378528 326898 378570 327134
rect 378806 326898 378848 327134
rect 378528 326866 378848 326898
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 378528 291454 378848 291486
rect 378528 291218 378570 291454
rect 378806 291218 378848 291454
rect 378528 291134 378848 291218
rect 378528 290898 378570 291134
rect 378806 290898 378848 291134
rect 378528 290866 378848 290898
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 378528 255454 378848 255486
rect 378528 255218 378570 255454
rect 378806 255218 378848 255454
rect 378528 255134 378848 255218
rect 378528 254898 378570 255134
rect 378806 254898 378848 255134
rect 378528 254866 378848 254898
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 389219 449716 389285 449717
rect 389219 449652 389220 449716
rect 389284 449652 389285 449716
rect 389219 449651 389285 449652
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 389222 109037 389282 449651
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 389219 109036 389285 109037
rect 389219 108972 389220 109036
rect 389284 108972 389285 109036
rect 389219 108971 389285 108972
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 415899 700500 415965 700501
rect 415899 700436 415900 700500
rect 415964 700436 415965 700500
rect 415899 700435 415965 700436
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 415902 457469 415962 700435
rect 416394 670054 417014 709082
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 418659 700364 418725 700365
rect 418659 700300 418660 700364
rect 418724 700300 418725 700364
rect 418659 700299 418725 700300
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 417923 622844 417989 622845
rect 417923 622780 417924 622844
rect 417988 622780 417989 622844
rect 417923 622779 417989 622780
rect 417555 618220 417621 618221
rect 417555 618156 417556 618220
rect 417620 618156 417621 618220
rect 417555 618155 417621 618156
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 417371 586940 417437 586941
rect 417371 586876 417372 586940
rect 417436 586876 417437 586940
rect 417371 586875 417437 586876
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 417374 494053 417434 586875
rect 417558 528189 417618 618155
rect 417739 586804 417805 586805
rect 417739 586740 417740 586804
rect 417804 586740 417805 586804
rect 417739 586739 417805 586740
rect 417555 528188 417621 528189
rect 417555 528124 417556 528188
rect 417620 528124 417621 528188
rect 417555 528123 417621 528124
rect 417558 527237 417618 528123
rect 417555 527236 417621 527237
rect 417555 527172 417556 527236
rect 417620 527172 417621 527236
rect 417555 527171 417621 527172
rect 417742 498133 417802 586739
rect 417926 532949 417986 622779
rect 417923 532948 417989 532949
rect 417923 532884 417924 532948
rect 417988 532884 417989 532948
rect 417923 532883 417989 532884
rect 417739 498132 417805 498133
rect 417739 498068 417740 498132
rect 417804 498068 417805 498132
rect 417739 498067 417805 498068
rect 417371 494052 417437 494053
rect 417371 493988 417372 494052
rect 417436 493988 417437 494052
rect 417371 493987 417437 493988
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 415899 457468 415965 457469
rect 415899 457404 415900 457468
rect 415964 457404 415965 457468
rect 415899 457403 415965 457404
rect 414611 454340 414677 454341
rect 414611 454276 414612 454340
rect 414676 454276 414677 454340
rect 414611 454275 414677 454276
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412674 306334 413294 341778
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 414614 17101 414674 454275
rect 416394 454054 417014 489498
rect 418662 480861 418722 700299
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 675244 424454 676938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 675244 434414 686898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 675244 438134 690618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 675244 441854 694338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 675244 445574 698058
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 675244 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 675244 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 675244 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 675244 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 675244 481574 698058
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 675244 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 675244 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 675244 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 675244 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 675244 517574 698058
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 675244 532454 676938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 675244 542414 686898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 675244 546134 690618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 675244 549854 694338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 675244 553574 698058
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 550955 674932 551021 674933
rect 550955 674868 550956 674932
rect 551020 674868 551021 674932
rect 550955 674867 551021 674868
rect 550958 673470 551018 674867
rect 550840 673410 551018 673470
rect 550840 673202 550900 673410
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 420272 655174 420620 655206
rect 420272 654938 420328 655174
rect 420564 654938 420620 655174
rect 420272 654854 420620 654938
rect 420272 654618 420328 654854
rect 420564 654618 420620 654854
rect 420272 654586 420620 654618
rect 556000 655174 556348 655206
rect 556000 654938 556056 655174
rect 556292 654938 556348 655174
rect 556000 654854 556348 654938
rect 556000 654618 556056 654854
rect 556292 654618 556348 654854
rect 556000 654586 556348 654618
rect 420952 651454 421300 651486
rect 420952 651218 421008 651454
rect 421244 651218 421300 651454
rect 420952 651134 421300 651218
rect 420952 650898 421008 651134
rect 421244 650898 421300 651134
rect 420952 650866 421300 650898
rect 555320 651454 555668 651486
rect 555320 651218 555376 651454
rect 555612 651218 555668 651454
rect 555320 651134 555668 651218
rect 555320 650898 555376 651134
rect 555612 650898 555668 651134
rect 555320 650866 555668 650898
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 420272 619174 420620 619206
rect 420272 618938 420328 619174
rect 420564 618938 420620 619174
rect 420272 618854 420620 618938
rect 420272 618618 420328 618854
rect 420564 618618 420620 618854
rect 420272 618586 420620 618618
rect 556000 619174 556348 619206
rect 556000 618938 556056 619174
rect 556292 618938 556348 619174
rect 556000 618854 556348 618938
rect 556000 618618 556056 618854
rect 556292 618618 556348 618854
rect 556000 618586 556348 618618
rect 420952 615454 421300 615486
rect 420952 615218 421008 615454
rect 421244 615218 421300 615454
rect 420952 615134 421300 615218
rect 420952 614898 421008 615134
rect 421244 614898 421300 615134
rect 420952 614866 421300 614898
rect 555320 615454 555668 615486
rect 555320 615218 555376 615454
rect 555612 615218 555668 615454
rect 555320 615134 555668 615218
rect 555320 614898 555376 615134
rect 555612 614898 555668 615134
rect 555320 614866 555668 614898
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 436056 589930 436116 590106
rect 437144 589930 437204 590106
rect 438232 589930 438292 590106
rect 436056 589870 436202 589930
rect 418843 587756 418909 587757
rect 418843 587692 418844 587756
rect 418908 587692 418909 587756
rect 418843 587691 418909 587692
rect 418846 493373 418906 587691
rect 436142 587077 436202 589870
rect 437062 589870 437204 589930
rect 438166 589870 438292 589930
rect 439592 589930 439652 590106
rect 440544 589930 440604 590106
rect 441768 589930 441828 590106
rect 439592 589870 439698 589930
rect 440544 589870 440618 589930
rect 437062 587893 437122 589870
rect 438166 587893 438226 589870
rect 439638 587893 439698 589870
rect 437059 587892 437125 587893
rect 437059 587828 437060 587892
rect 437124 587828 437125 587892
rect 437059 587827 437125 587828
rect 438163 587892 438229 587893
rect 438163 587828 438164 587892
rect 438228 587828 438229 587892
rect 438163 587827 438229 587828
rect 439635 587892 439701 587893
rect 439635 587828 439636 587892
rect 439700 587828 439701 587892
rect 439635 587827 439701 587828
rect 419763 587076 419829 587077
rect 419763 587012 419764 587076
rect 419828 587012 419829 587076
rect 419763 587011 419829 587012
rect 436139 587076 436205 587077
rect 436139 587012 436140 587076
rect 436204 587012 436205 587076
rect 436139 587011 436205 587012
rect 419395 584900 419461 584901
rect 419395 584836 419396 584900
rect 419460 584836 419461 584900
rect 419395 584835 419461 584836
rect 419398 497997 419458 584835
rect 419395 497996 419461 497997
rect 419395 497932 419396 497996
rect 419460 497932 419461 497996
rect 419395 497931 419461 497932
rect 419766 496773 419826 587011
rect 440558 586805 440618 589870
rect 441662 589870 441828 589930
rect 443128 589930 443188 590106
rect 444216 589930 444276 590106
rect 445440 589930 445500 590106
rect 446528 589930 446588 590106
rect 447616 589930 447676 590106
rect 448296 589930 448356 590106
rect 448704 589930 448764 590106
rect 450064 589930 450124 590106
rect 450744 589930 450804 590106
rect 451288 589930 451348 590106
rect 452376 589930 452436 590106
rect 453464 589930 453524 590106
rect 443128 589870 443194 589930
rect 444216 589870 444298 589930
rect 445440 589870 445586 589930
rect 441662 587893 441722 589870
rect 443134 587893 443194 589870
rect 444238 587893 444298 589870
rect 445526 587893 445586 589870
rect 446446 589870 446588 589930
rect 447550 589870 447676 589930
rect 448286 589870 448356 589930
rect 448654 589870 448764 589930
rect 449942 589870 450124 589930
rect 450678 589870 450804 589930
rect 451046 589870 451348 589930
rect 452334 589870 452436 589930
rect 453438 589870 453524 589930
rect 453600 589930 453660 590106
rect 454552 589930 454612 590106
rect 455912 589930 455972 590106
rect 453600 589870 453682 589930
rect 446446 587893 446506 589870
rect 447550 587893 447610 589870
rect 441659 587892 441725 587893
rect 441659 587828 441660 587892
rect 441724 587828 441725 587892
rect 441659 587827 441725 587828
rect 443131 587892 443197 587893
rect 443131 587828 443132 587892
rect 443196 587828 443197 587892
rect 443131 587827 443197 587828
rect 444235 587892 444301 587893
rect 444235 587828 444236 587892
rect 444300 587828 444301 587892
rect 444235 587827 444301 587828
rect 445523 587892 445589 587893
rect 445523 587828 445524 587892
rect 445588 587828 445589 587892
rect 445523 587827 445589 587828
rect 446443 587892 446509 587893
rect 446443 587828 446444 587892
rect 446508 587828 446509 587892
rect 446443 587827 446509 587828
rect 447547 587892 447613 587893
rect 447547 587828 447548 587892
rect 447612 587828 447613 587892
rect 447547 587827 447613 587828
rect 448286 587757 448346 589870
rect 448654 587893 448714 589870
rect 449942 587893 450002 589870
rect 450678 587893 450738 589870
rect 448651 587892 448717 587893
rect 448651 587828 448652 587892
rect 448716 587828 448717 587892
rect 448651 587827 448717 587828
rect 449939 587892 450005 587893
rect 449939 587828 449940 587892
rect 450004 587828 450005 587892
rect 449939 587827 450005 587828
rect 450675 587892 450741 587893
rect 450675 587828 450676 587892
rect 450740 587828 450741 587892
rect 450675 587827 450741 587828
rect 448283 587756 448349 587757
rect 448283 587692 448284 587756
rect 448348 587692 448349 587756
rect 448283 587691 448349 587692
rect 451046 587210 451106 589870
rect 452334 587757 452394 589870
rect 453438 587757 453498 589870
rect 453622 587893 453682 589870
rect 454542 589870 454612 589930
rect 455830 589870 455972 589930
rect 456048 589930 456108 590106
rect 457000 589930 457060 590106
rect 458088 589930 458148 590106
rect 458496 589930 458556 590106
rect 459448 589930 459508 590106
rect 460672 589930 460732 590106
rect 461080 589930 461140 590106
rect 461760 589930 461820 590106
rect 462848 589930 462908 590106
rect 456048 589870 456258 589930
rect 454542 587893 454602 589870
rect 453619 587892 453685 587893
rect 453619 587828 453620 587892
rect 453684 587828 453685 587892
rect 453619 587827 453685 587828
rect 454539 587892 454605 587893
rect 454539 587828 454540 587892
rect 454604 587828 454605 587892
rect 454539 587827 454605 587828
rect 455830 587757 455890 589870
rect 456198 587893 456258 589870
rect 456934 589870 457060 589930
rect 458038 589870 458148 589930
rect 458406 589870 458556 589930
rect 459326 589870 459508 589930
rect 460614 589870 460732 589930
rect 460982 589870 461140 589930
rect 461718 589870 461820 589930
rect 462822 589870 462908 589930
rect 463528 589930 463588 590106
rect 463936 589930 463996 590106
rect 465296 589930 465356 590106
rect 465976 589930 466036 590106
rect 466384 589930 466444 590106
rect 467608 589930 467668 590106
rect 463528 589870 463618 589930
rect 456934 587893 456994 589870
rect 458038 587893 458098 589870
rect 456195 587892 456261 587893
rect 456195 587828 456196 587892
rect 456260 587828 456261 587892
rect 456195 587827 456261 587828
rect 456931 587892 456997 587893
rect 456931 587828 456932 587892
rect 456996 587828 456997 587892
rect 456931 587827 456997 587828
rect 458035 587892 458101 587893
rect 458035 587828 458036 587892
rect 458100 587828 458101 587892
rect 458035 587827 458101 587828
rect 452331 587756 452397 587757
rect 452331 587692 452332 587756
rect 452396 587692 452397 587756
rect 452331 587691 452397 587692
rect 453435 587756 453501 587757
rect 453435 587692 453436 587756
rect 453500 587692 453501 587756
rect 453435 587691 453501 587692
rect 455827 587756 455893 587757
rect 455827 587692 455828 587756
rect 455892 587692 455893 587756
rect 455827 587691 455893 587692
rect 458406 587213 458466 589870
rect 459326 587757 459386 589870
rect 460614 587757 460674 589870
rect 460982 587757 461042 589870
rect 461718 587757 461778 589870
rect 459323 587756 459389 587757
rect 459323 587692 459324 587756
rect 459388 587692 459389 587756
rect 459323 587691 459389 587692
rect 460611 587756 460677 587757
rect 460611 587692 460612 587756
rect 460676 587692 460677 587756
rect 460611 587691 460677 587692
rect 460979 587756 461045 587757
rect 460979 587692 460980 587756
rect 461044 587692 461045 587756
rect 460979 587691 461045 587692
rect 461715 587756 461781 587757
rect 461715 587692 461716 587756
rect 461780 587692 461781 587756
rect 461715 587691 461781 587692
rect 462822 587213 462882 589870
rect 463558 587757 463618 589870
rect 463926 589870 463996 589930
rect 465214 589870 465356 589930
rect 465950 589870 466036 589930
rect 466318 589870 466444 589930
rect 467606 589870 467668 589930
rect 468288 589930 468348 590106
rect 468696 589930 468756 590106
rect 469784 589930 469844 590106
rect 471008 589930 471068 590106
rect 468288 589870 468402 589930
rect 468696 589870 468770 589930
rect 469784 589870 469874 589930
rect 463926 587757 463986 589870
rect 463555 587756 463621 587757
rect 463555 587692 463556 587756
rect 463620 587692 463621 587756
rect 463555 587691 463621 587692
rect 463923 587756 463989 587757
rect 463923 587692 463924 587756
rect 463988 587692 463989 587756
rect 463923 587691 463989 587692
rect 465214 587213 465274 589870
rect 465950 587757 466010 589870
rect 466318 587757 466378 589870
rect 467606 587757 467666 589870
rect 465947 587756 466013 587757
rect 465947 587692 465948 587756
rect 466012 587692 466013 587756
rect 465947 587691 466013 587692
rect 466315 587756 466381 587757
rect 466315 587692 466316 587756
rect 466380 587692 466381 587756
rect 466315 587691 466381 587692
rect 467603 587756 467669 587757
rect 467603 587692 467604 587756
rect 467668 587692 467669 587756
rect 467603 587691 467669 587692
rect 458403 587212 458469 587213
rect 451046 587150 451474 587210
rect 451414 586941 451474 587150
rect 458403 587148 458404 587212
rect 458468 587148 458469 587212
rect 458403 587147 458469 587148
rect 462819 587212 462885 587213
rect 462819 587148 462820 587212
rect 462884 587148 462885 587212
rect 462819 587147 462885 587148
rect 465211 587212 465277 587213
rect 465211 587148 465212 587212
rect 465276 587148 465277 587212
rect 465211 587147 465277 587148
rect 468342 587077 468402 589870
rect 468710 587757 468770 589870
rect 469814 587757 469874 589870
rect 470366 589870 471068 589930
rect 471144 589930 471204 590106
rect 472232 589930 472292 590106
rect 473320 589930 473380 590106
rect 473592 589930 473652 590106
rect 471144 589870 471346 589930
rect 468707 587756 468773 587757
rect 468707 587692 468708 587756
rect 468772 587692 468773 587756
rect 468707 587691 468773 587692
rect 469811 587756 469877 587757
rect 469811 587692 469812 587756
rect 469876 587692 469877 587756
rect 469811 587691 469877 587692
rect 468339 587076 468405 587077
rect 468339 587012 468340 587076
rect 468404 587012 468405 587076
rect 468339 587011 468405 587012
rect 451411 586940 451477 586941
rect 451411 586876 451412 586940
rect 451476 586876 451477 586940
rect 451411 586875 451477 586876
rect 440555 586804 440621 586805
rect 440555 586740 440556 586804
rect 440620 586740 440621 586804
rect 440555 586739 440621 586740
rect 470366 586530 470426 589870
rect 471286 587893 471346 589870
rect 472206 589870 472292 589930
rect 473310 589870 473380 589930
rect 473494 589870 473652 589930
rect 474408 589930 474468 590106
rect 475768 589930 475828 590106
rect 474408 589870 474474 589930
rect 472206 587893 472266 589870
rect 473310 587893 473370 589870
rect 471283 587892 471349 587893
rect 471283 587828 471284 587892
rect 471348 587828 471349 587892
rect 471283 587827 471349 587828
rect 472203 587892 472269 587893
rect 472203 587828 472204 587892
rect 472268 587828 472269 587892
rect 472203 587827 472269 587828
rect 473307 587892 473373 587893
rect 473307 587828 473308 587892
rect 473372 587828 473373 587892
rect 473307 587827 473373 587828
rect 473494 587621 473554 589870
rect 474414 587893 474474 589870
rect 475702 589870 475828 589930
rect 476040 589930 476100 590106
rect 476992 589930 477052 590106
rect 476040 589870 476130 589930
rect 474411 587892 474477 587893
rect 474411 587828 474412 587892
rect 474476 587828 474477 587892
rect 474411 587827 474477 587828
rect 473491 587620 473557 587621
rect 473491 587556 473492 587620
rect 473556 587556 473557 587620
rect 473491 587555 473557 587556
rect 475702 586941 475762 589870
rect 476070 587485 476130 589870
rect 476990 589870 477052 589930
rect 478080 589930 478140 590106
rect 478488 589930 478548 590106
rect 478080 589870 478154 589930
rect 476990 587893 477050 589870
rect 478094 587893 478154 589870
rect 478462 589870 478548 589930
rect 479168 589930 479228 590106
rect 480936 589930 480996 590106
rect 483520 589930 483580 590106
rect 479168 589870 479258 589930
rect 476987 587892 477053 587893
rect 476987 587828 476988 587892
rect 477052 587828 477053 587892
rect 476987 587827 477053 587828
rect 478091 587892 478157 587893
rect 478091 587828 478092 587892
rect 478156 587828 478157 587892
rect 478091 587827 478157 587828
rect 476067 587484 476133 587485
rect 476067 587420 476068 587484
rect 476132 587420 476133 587484
rect 476067 587419 476133 587420
rect 478462 587349 478522 589870
rect 479198 587893 479258 589870
rect 480854 589870 480996 589930
rect 483430 589870 483580 589930
rect 485968 589930 486028 590106
rect 488280 589930 488340 590106
rect 491000 589930 491060 590106
rect 493448 589930 493508 590106
rect 485968 589870 486066 589930
rect 480854 587893 480914 589870
rect 483430 587893 483490 589870
rect 486006 587893 486066 589870
rect 488214 589870 488340 589930
rect 490974 589870 491060 589930
rect 493366 589870 493508 589930
rect 495896 589930 495956 590106
rect 498480 589930 498540 590106
rect 500928 589930 500988 590106
rect 503512 589930 503572 590106
rect 505960 589930 506020 590106
rect 508544 589930 508604 590106
rect 495896 589870 496002 589930
rect 498480 589870 498578 589930
rect 488214 587893 488274 589870
rect 490974 589290 491034 589870
rect 489686 589230 491034 589290
rect 479195 587892 479261 587893
rect 479195 587828 479196 587892
rect 479260 587828 479261 587892
rect 479195 587827 479261 587828
rect 480851 587892 480917 587893
rect 480851 587828 480852 587892
rect 480916 587828 480917 587892
rect 480851 587827 480917 587828
rect 483427 587892 483493 587893
rect 483427 587828 483428 587892
rect 483492 587828 483493 587892
rect 483427 587827 483493 587828
rect 486003 587892 486069 587893
rect 486003 587828 486004 587892
rect 486068 587828 486069 587892
rect 486003 587827 486069 587828
rect 488211 587892 488277 587893
rect 488211 587828 488212 587892
rect 488276 587828 488277 587892
rect 488211 587827 488277 587828
rect 478459 587348 478525 587349
rect 478459 587284 478460 587348
rect 478524 587284 478525 587348
rect 478459 587283 478525 587284
rect 475699 586940 475765 586941
rect 475699 586876 475700 586940
rect 475764 586876 475765 586940
rect 475699 586875 475765 586876
rect 470547 586532 470613 586533
rect 470547 586530 470548 586532
rect 470366 586470 470548 586530
rect 470547 586468 470548 586470
rect 470612 586468 470613 586532
rect 489686 586530 489746 589230
rect 493366 587893 493426 589870
rect 495942 587893 496002 589870
rect 498518 587893 498578 589870
rect 500910 589870 500988 589930
rect 503486 589870 503572 589930
rect 505878 589870 506020 589930
rect 508454 589870 508604 589930
rect 510992 589930 511052 590106
rect 513440 589930 513500 590106
rect 515888 589930 515948 590106
rect 518472 589930 518532 590106
rect 510992 589870 511090 589930
rect 500910 587893 500970 589870
rect 503486 587893 503546 589870
rect 505878 587893 505938 589870
rect 508454 587893 508514 589870
rect 511030 587893 511090 589870
rect 513422 589870 513500 589930
rect 515814 589870 515948 589930
rect 518390 589870 518532 589930
rect 520920 589930 520980 590106
rect 523368 589930 523428 590106
rect 525952 589930 526012 590106
rect 520920 589870 521026 589930
rect 513422 587893 513482 589870
rect 515814 587893 515874 589870
rect 518390 587893 518450 589870
rect 520966 587893 521026 589870
rect 523358 589870 523428 589930
rect 525934 589870 526012 589930
rect 523358 587893 523418 589870
rect 525934 587893 525994 589870
rect 493363 587892 493429 587893
rect 493363 587828 493364 587892
rect 493428 587828 493429 587892
rect 493363 587827 493429 587828
rect 495939 587892 496005 587893
rect 495939 587828 495940 587892
rect 496004 587828 496005 587892
rect 495939 587827 496005 587828
rect 498515 587892 498581 587893
rect 498515 587828 498516 587892
rect 498580 587828 498581 587892
rect 498515 587827 498581 587828
rect 500907 587892 500973 587893
rect 500907 587828 500908 587892
rect 500972 587828 500973 587892
rect 500907 587827 500973 587828
rect 503483 587892 503549 587893
rect 503483 587828 503484 587892
rect 503548 587828 503549 587892
rect 503483 587827 503549 587828
rect 505875 587892 505941 587893
rect 505875 587828 505876 587892
rect 505940 587828 505941 587892
rect 505875 587827 505941 587828
rect 508451 587892 508517 587893
rect 508451 587828 508452 587892
rect 508516 587828 508517 587892
rect 508451 587827 508517 587828
rect 511027 587892 511093 587893
rect 511027 587828 511028 587892
rect 511092 587828 511093 587892
rect 511027 587827 511093 587828
rect 513419 587892 513485 587893
rect 513419 587828 513420 587892
rect 513484 587828 513485 587892
rect 513419 587827 513485 587828
rect 515811 587892 515877 587893
rect 515811 587828 515812 587892
rect 515876 587828 515877 587892
rect 515811 587827 515877 587828
rect 517467 587892 517533 587893
rect 517467 587828 517468 587892
rect 517532 587828 517533 587892
rect 517467 587827 517533 587828
rect 518387 587892 518453 587893
rect 518387 587828 518388 587892
rect 518452 587828 518453 587892
rect 518387 587827 518453 587828
rect 520963 587892 521029 587893
rect 520963 587828 520964 587892
rect 521028 587828 521029 587892
rect 520963 587827 521029 587828
rect 523355 587892 523421 587893
rect 523355 587828 523356 587892
rect 523420 587828 523421 587892
rect 523355 587827 523421 587828
rect 525931 587892 525997 587893
rect 525931 587828 525932 587892
rect 525996 587828 525997 587892
rect 525931 587827 525997 587828
rect 489867 586532 489933 586533
rect 489867 586530 489868 586532
rect 489686 586470 489868 586530
rect 470547 586467 470613 586468
rect 489867 586468 489868 586470
rect 489932 586468 489933 586532
rect 489867 586467 489933 586468
rect 517470 585717 517530 587827
rect 517467 585716 517533 585717
rect 517467 585652 517468 585716
rect 517532 585652 517533 585716
rect 517467 585651 517533 585652
rect 550771 585308 550837 585309
rect 550771 585244 550772 585308
rect 550836 585244 550837 585308
rect 550771 585243 550837 585244
rect 550774 583810 550834 585243
rect 550774 583750 550900 583810
rect 550840 583202 550900 583750
rect 420272 582929 420620 583036
rect 420272 582693 420328 582929
rect 420564 582693 420620 582929
rect 420272 582586 420620 582693
rect 556000 582929 556348 583036
rect 556000 582693 556056 582929
rect 556292 582693 556348 582929
rect 556000 582586 556348 582693
rect 420952 579454 421300 579486
rect 420952 579218 421008 579454
rect 421244 579218 421300 579454
rect 420952 579134 421300 579218
rect 420952 578898 421008 579134
rect 421244 578898 421300 579134
rect 420952 578866 421300 578898
rect 555320 579454 555668 579486
rect 555320 579218 555376 579454
rect 555612 579218 555668 579454
rect 555320 579134 555668 579218
rect 555320 578898 555376 579134
rect 555612 578898 555668 579134
rect 555320 578866 555668 578898
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 420272 547174 420620 547206
rect 420272 546938 420328 547174
rect 420564 546938 420620 547174
rect 420272 546854 420620 546938
rect 420272 546618 420328 546854
rect 420564 546618 420620 546854
rect 420272 546586 420620 546618
rect 556000 547174 556348 547206
rect 556000 546938 556056 547174
rect 556292 546938 556348 547174
rect 556000 546854 556348 546938
rect 556000 546618 556056 546854
rect 556292 546618 556348 546854
rect 556000 546586 556348 546618
rect 420952 543454 421300 543486
rect 420952 543218 421008 543454
rect 421244 543218 421300 543454
rect 420952 543134 421300 543218
rect 420952 542898 421008 543134
rect 421244 542898 421300 543134
rect 420952 542866 421300 542898
rect 555320 543454 555668 543486
rect 555320 543218 555376 543454
rect 555612 543218 555668 543454
rect 555320 543134 555668 543218
rect 555320 542898 555376 543134
rect 555612 542898 555668 543134
rect 555320 542866 555668 542898
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 420272 511174 420620 511206
rect 420272 510938 420328 511174
rect 420564 510938 420620 511174
rect 420272 510854 420620 510938
rect 420272 510618 420328 510854
rect 420564 510618 420620 510854
rect 420272 510586 420620 510618
rect 556000 511174 556348 511206
rect 556000 510938 556056 511174
rect 556292 510938 556348 511174
rect 556000 510854 556348 510938
rect 556000 510618 556056 510854
rect 556292 510618 556348 510854
rect 556000 510586 556348 510618
rect 420952 507454 421300 507486
rect 420952 507218 421008 507454
rect 421244 507218 421300 507454
rect 420952 507134 421300 507218
rect 420952 506898 421008 507134
rect 421244 506898 421300 507134
rect 420952 506866 421300 506898
rect 555320 507454 555668 507486
rect 555320 507218 555376 507454
rect 555612 507218 555668 507454
rect 555320 507134 555668 507218
rect 555320 506898 555376 507134
rect 555612 506898 555668 507134
rect 555320 506866 555668 506898
rect 436056 499590 436116 500106
rect 437144 499590 437204 500106
rect 436056 499530 436202 499590
rect 419763 496772 419829 496773
rect 419763 496708 419764 496772
rect 419828 496708 419829 496772
rect 419763 496707 419829 496708
rect 420114 493774 420734 498064
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 418843 493372 418909 493373
rect 418843 493308 418844 493372
rect 418908 493308 418909 493372
rect 418843 493307 418909 493308
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 418659 480860 418725 480861
rect 418659 480796 418660 480860
rect 418724 480796 418725 480860
rect 418659 480795 418725 480796
rect 417371 463724 417437 463725
rect 417371 463660 417372 463724
rect 417436 463660 417437 463724
rect 417371 463659 417437 463660
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 415899 451892 415965 451893
rect 415899 451828 415900 451892
rect 415964 451828 415965 451892
rect 415899 451827 415965 451828
rect 415902 19277 415962 451827
rect 416083 449852 416149 449853
rect 416083 449788 416084 449852
rect 416148 449788 416149 449852
rect 416083 449787 416149 449788
rect 415899 19276 415965 19277
rect 415899 19212 415900 19276
rect 415964 19212 415965 19276
rect 415899 19211 415965 19212
rect 414611 17100 414677 17101
rect 414611 17036 414612 17100
rect 414676 17036 414677 17100
rect 414611 17035 414677 17036
rect 416086 16693 416146 449787
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 416394 310054 417014 345498
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 130054 417014 165498
rect 417187 146028 417253 146029
rect 417187 145964 417188 146028
rect 417252 145964 417253 146028
rect 417187 145963 417253 145964
rect 416394 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 417014 130054
rect 416394 129734 417014 129818
rect 416394 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 417014 129734
rect 416394 94054 417014 129498
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 417190 55997 417250 145963
rect 417374 107541 417434 463659
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 418107 453116 418173 453117
rect 418107 453052 418108 453116
rect 418172 453052 418173 453116
rect 418107 453051 418173 453052
rect 417739 450940 417805 450941
rect 417739 450876 417740 450940
rect 417804 450876 417805 450940
rect 417739 450875 417805 450876
rect 417555 449172 417621 449173
rect 417555 449108 417556 449172
rect 417620 449108 417621 449172
rect 417555 449107 417621 449108
rect 417558 138277 417618 449107
rect 417742 146029 417802 450875
rect 417739 146028 417805 146029
rect 417739 145964 417740 146028
rect 417804 145964 417805 146028
rect 417739 145963 417805 145964
rect 417739 142764 417805 142765
rect 417739 142700 417740 142764
rect 417804 142700 417805 142764
rect 417739 142699 417805 142700
rect 417555 138276 417621 138277
rect 417555 138212 417556 138276
rect 417620 138212 417621 138276
rect 417555 138211 417621 138212
rect 417371 107540 417437 107541
rect 417371 107476 417372 107540
rect 417436 107476 417437 107540
rect 417371 107475 417437 107476
rect 417187 55996 417253 55997
rect 417187 55932 417188 55996
rect 417252 55932 417253 55996
rect 417187 55931 417253 55932
rect 417742 52869 417802 142699
rect 417923 138276 417989 138277
rect 417923 138212 417924 138276
rect 417988 138212 417989 138276
rect 417923 138211 417989 138212
rect 417739 52868 417805 52869
rect 417739 52804 417740 52868
rect 417804 52804 417805 52868
rect 417739 52803 417805 52804
rect 417926 48245 417986 138211
rect 417923 48244 417989 48245
rect 417923 48180 417924 48244
rect 417988 48180 417989 48244
rect 417923 48179 417989 48180
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416083 16692 416149 16693
rect 416083 16628 416084 16692
rect 416148 16628 416149 16692
rect 416083 16627 416149 16628
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 -5146 417014 21498
rect 418110 19141 418170 453051
rect 418659 452436 418725 452437
rect 418659 452372 418660 452436
rect 418724 452372 418725 452436
rect 418659 452371 418725 452372
rect 418107 19140 418173 19141
rect 418107 19076 418108 19140
rect 418172 19076 418173 19140
rect 418107 19075 418173 19076
rect 418662 19005 418722 452371
rect 418843 452300 418909 452301
rect 418843 452236 418844 452300
rect 418908 452236 418909 452300
rect 418843 452235 418909 452236
rect 418846 19141 418906 452235
rect 419027 451756 419093 451757
rect 419027 451692 419028 451756
rect 419092 451692 419093 451756
rect 419027 451691 419093 451692
rect 419030 106997 419090 451691
rect 420114 421774 420734 457218
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 420114 313774 420734 349218
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 195244 420734 205218
rect 423834 497494 424454 498064
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 425494 424454 460938
rect 423834 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 424454 425494
rect 423834 425174 424454 425258
rect 423834 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 424454 425174
rect 423834 389494 424454 424938
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 423834 317494 424454 352938
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 195244 424454 208938
rect 433794 471454 434414 498064
rect 436142 496909 436202 499530
rect 437062 499530 437204 499590
rect 438232 499590 438292 500106
rect 439592 499590 439652 500106
rect 440544 499590 440604 500106
rect 441768 499590 441828 500106
rect 438232 499530 438410 499590
rect 439592 499530 439698 499590
rect 440544 499530 440618 499590
rect 437062 497045 437122 499530
rect 437059 497044 437125 497045
rect 437059 496980 437060 497044
rect 437124 496980 437125 497044
rect 437059 496979 437125 496980
rect 436139 496908 436205 496909
rect 436139 496844 436140 496908
rect 436204 496844 436205 496908
rect 436139 496843 436205 496844
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 195244 434414 218898
rect 437514 475174 438134 498064
rect 438350 496909 438410 499530
rect 439638 496909 439698 499530
rect 440558 498133 440618 499530
rect 441662 499530 441828 499590
rect 443128 499590 443188 500106
rect 444216 499590 444276 500106
rect 445440 499590 445500 500106
rect 443128 499530 443194 499590
rect 444216 499530 444298 499590
rect 441662 498133 441722 499530
rect 440555 498132 440621 498133
rect 440555 498068 440556 498132
rect 440620 498068 440621 498132
rect 440555 498067 440621 498068
rect 441659 498132 441725 498133
rect 441659 498068 441660 498132
rect 441724 498068 441725 498132
rect 441659 498067 441725 498068
rect 440558 496909 440618 498067
rect 438347 496908 438413 496909
rect 438347 496844 438348 496908
rect 438412 496844 438413 496908
rect 438347 496843 438413 496844
rect 439635 496908 439701 496909
rect 439635 496844 439636 496908
rect 439700 496844 439701 496908
rect 439635 496843 439701 496844
rect 440555 496908 440621 496909
rect 440555 496844 440556 496908
rect 440620 496844 440621 496908
rect 440555 496843 440621 496844
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 195244 438134 222618
rect 441234 478894 441854 497940
rect 443134 496909 443194 499530
rect 444238 497453 444298 499530
rect 445342 499530 445500 499590
rect 446528 499590 446588 500106
rect 447616 499590 447676 500106
rect 448296 499590 448356 500106
rect 448704 499590 448764 500106
rect 446528 499530 446690 499590
rect 447616 499530 447794 499590
rect 445342 498133 445402 499530
rect 445339 498132 445405 498133
rect 445339 498068 445340 498132
rect 445404 498068 445405 498132
rect 445339 498067 445405 498068
rect 444235 497452 444301 497453
rect 444235 497388 444236 497452
rect 444300 497388 444301 497452
rect 444235 497387 444301 497388
rect 443131 496908 443197 496909
rect 443131 496844 443132 496908
rect 443196 496844 443197 496908
rect 443131 496843 443197 496844
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 195244 441854 226338
rect 444954 482614 445574 497940
rect 446630 497181 446690 499530
rect 446627 497180 446693 497181
rect 446627 497116 446628 497180
rect 446692 497116 446693 497180
rect 446627 497115 446693 497116
rect 447734 497045 447794 499530
rect 448286 499530 448356 499590
rect 448654 499530 448764 499590
rect 450064 499590 450124 500106
rect 450744 499590 450804 500106
rect 450064 499530 450186 499590
rect 447731 497044 447797 497045
rect 447731 496980 447732 497044
rect 447796 496980 447797 497044
rect 447731 496979 447797 496980
rect 448286 496909 448346 499530
rect 448654 498133 448714 499530
rect 448651 498132 448717 498133
rect 448651 498068 448652 498132
rect 448716 498068 448717 498132
rect 448651 498067 448717 498068
rect 448283 496908 448349 496909
rect 448283 496844 448284 496908
rect 448348 496844 448349 496908
rect 448283 496843 448349 496844
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 195244 445574 230058
rect 448674 486334 449294 497940
rect 450126 497453 450186 499530
rect 450678 499530 450804 499590
rect 450123 497452 450189 497453
rect 450123 497388 450124 497452
rect 450188 497388 450189 497452
rect 450123 497387 450189 497388
rect 450678 496909 450738 499530
rect 451288 499490 451348 500106
rect 452376 499590 452436 500106
rect 453464 499590 453524 500106
rect 451046 499430 451348 499490
rect 452334 499530 452436 499590
rect 453438 499530 453524 499590
rect 453600 499590 453660 500106
rect 454552 499590 454612 500106
rect 455912 499590 455972 500106
rect 453600 499530 453682 499590
rect 451046 498133 451106 499430
rect 452334 498133 452394 499530
rect 451043 498132 451109 498133
rect 451043 498068 451044 498132
rect 451108 498068 451109 498132
rect 451043 498067 451109 498068
rect 452331 498132 452397 498133
rect 452331 498068 452332 498132
rect 452396 498068 452397 498132
rect 452331 498067 452397 498068
rect 450675 496908 450741 496909
rect 450675 496844 450676 496908
rect 450740 496844 450741 496908
rect 450675 496843 450741 496844
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448674 306334 449294 341778
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 195244 449294 197778
rect 452394 490054 453014 497940
rect 453438 497045 453498 499530
rect 453435 497044 453501 497045
rect 453435 496980 453436 497044
rect 453500 496980 453501 497044
rect 453435 496979 453501 496980
rect 453622 496909 453682 499530
rect 454542 499530 454612 499590
rect 455830 499530 455972 499590
rect 456048 499590 456108 500106
rect 457000 499590 457060 500106
rect 458088 499590 458148 500106
rect 458496 499590 458556 500106
rect 456048 499530 456258 499590
rect 454542 498133 454602 499530
rect 454539 498132 454605 498133
rect 454539 498068 454540 498132
rect 454604 498068 454605 498132
rect 454539 498067 454605 498068
rect 455830 496909 455890 499530
rect 456198 498133 456258 499530
rect 456934 499530 457060 499590
rect 458038 499530 458148 499590
rect 458406 499530 458556 499590
rect 459448 499590 459508 500106
rect 460672 499590 460732 500106
rect 461080 499590 461140 500106
rect 461760 499590 461820 500106
rect 462848 499590 462908 500106
rect 459448 499530 459570 499590
rect 456195 498132 456261 498133
rect 456195 498068 456196 498132
rect 456260 498068 456261 498132
rect 456195 498067 456261 498068
rect 453619 496908 453685 496909
rect 453619 496844 453620 496908
rect 453684 496844 453685 496908
rect 453619 496843 453685 496844
rect 455827 496908 455893 496909
rect 455827 496844 455828 496908
rect 455892 496844 455893 496908
rect 455827 496843 455893 496844
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 452394 310054 453014 345498
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 195244 453014 201498
rect 456114 493774 456734 497940
rect 456934 496909 456994 499530
rect 458038 497453 458098 499530
rect 458035 497452 458101 497453
rect 458035 497388 458036 497452
rect 458100 497388 458101 497452
rect 458035 497387 458101 497388
rect 458406 496909 458466 499530
rect 459510 496909 459570 499530
rect 460614 499530 460732 499590
rect 460982 499530 461140 499590
rect 461718 499530 461820 499590
rect 462822 499530 462908 499590
rect 463528 499590 463588 500106
rect 463936 499590 463996 500106
rect 465296 499590 465356 500106
rect 465976 499590 466036 500106
rect 466384 499590 466444 500106
rect 467608 499590 467668 500106
rect 463528 499530 463618 499590
rect 459834 497494 460454 498064
rect 460614 497861 460674 499530
rect 460611 497860 460677 497861
rect 460611 497796 460612 497860
rect 460676 497796 460677 497860
rect 460611 497795 460677 497796
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 456931 496908 456997 496909
rect 456931 496844 456932 496908
rect 456996 496844 456997 496908
rect 456931 496843 456997 496844
rect 458403 496908 458469 496909
rect 458403 496844 458404 496908
rect 458468 496844 458469 496908
rect 458403 496843 458469 496844
rect 459507 496908 459573 496909
rect 459507 496844 459508 496908
rect 459572 496844 459573 496908
rect 459507 496843 459573 496844
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 195244 456734 205218
rect 459834 461494 460454 496938
rect 460982 496909 461042 499530
rect 461718 497317 461778 499530
rect 462822 497861 462882 499530
rect 462819 497860 462885 497861
rect 462819 497796 462820 497860
rect 462884 497796 462885 497860
rect 462819 497795 462885 497796
rect 461715 497316 461781 497317
rect 461715 497252 461716 497316
rect 461780 497252 461781 497316
rect 461715 497251 461781 497252
rect 463558 496909 463618 499530
rect 463926 499530 463996 499590
rect 465214 499530 465356 499590
rect 465950 499530 466036 499590
rect 466318 499530 466444 499590
rect 467606 499530 467668 499590
rect 468288 499590 468348 500106
rect 468696 499590 468756 500106
rect 469784 499590 469844 500106
rect 471008 499590 471068 500106
rect 468288 499530 468402 499590
rect 468696 499530 468770 499590
rect 469784 499530 469874 499590
rect 463926 497997 463986 499530
rect 463923 497996 463989 497997
rect 463923 497932 463924 497996
rect 463988 497932 463989 497996
rect 463923 497931 463989 497932
rect 465214 497181 465274 499530
rect 465211 497180 465277 497181
rect 465211 497116 465212 497180
rect 465276 497116 465277 497180
rect 465211 497115 465277 497116
rect 465950 496909 466010 499530
rect 466318 497317 466378 499530
rect 467606 497453 467666 499530
rect 467603 497452 467669 497453
rect 467603 497388 467604 497452
rect 467668 497388 467669 497452
rect 467603 497387 467669 497388
rect 466315 497316 466381 497317
rect 466315 497252 466316 497316
rect 466380 497252 466381 497316
rect 466315 497251 466381 497252
rect 468342 496909 468402 499530
rect 468710 497997 468770 499530
rect 469814 498133 469874 499530
rect 470918 499530 471068 499590
rect 471144 499590 471204 500106
rect 472232 499590 472292 500106
rect 473320 499590 473380 500106
rect 471144 499530 471346 499590
rect 469811 498132 469877 498133
rect 469811 498068 469812 498132
rect 469876 498068 469877 498132
rect 469811 498067 469877 498068
rect 468707 497996 468773 497997
rect 468707 497932 468708 497996
rect 468772 497932 468773 497996
rect 468707 497931 468773 497932
rect 460979 496908 461045 496909
rect 460979 496844 460980 496908
rect 461044 496844 461045 496908
rect 460979 496843 461045 496844
rect 463555 496908 463621 496909
rect 463555 496844 463556 496908
rect 463620 496844 463621 496908
rect 463555 496843 463621 496844
rect 465947 496908 466013 496909
rect 465947 496844 465948 496908
rect 466012 496844 466013 496908
rect 465947 496843 466013 496844
rect 468339 496908 468405 496909
rect 468339 496844 468340 496908
rect 468404 496844 468405 496908
rect 468339 496843 468405 496844
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 195244 460454 208938
rect 469794 471454 470414 497940
rect 470918 496909 470978 499530
rect 471286 497725 471346 499530
rect 472206 499530 472292 499590
rect 473310 499530 473380 499590
rect 473592 499590 473652 500106
rect 474408 499590 474468 500106
rect 475768 499590 475828 500106
rect 473592 499530 473738 499590
rect 474408 499530 474474 499590
rect 471283 497724 471349 497725
rect 471283 497660 471284 497724
rect 471348 497660 471349 497724
rect 471283 497659 471349 497660
rect 472206 497045 472266 499530
rect 473310 498133 473370 499530
rect 473678 498133 473738 499530
rect 473307 498132 473373 498133
rect 473307 498068 473308 498132
rect 473372 498068 473373 498132
rect 473307 498067 473373 498068
rect 473675 498132 473741 498133
rect 473675 498068 473676 498132
rect 473740 498068 473741 498132
rect 473675 498067 473741 498068
rect 472203 497044 472269 497045
rect 472203 496980 472204 497044
rect 472268 496980 472269 497044
rect 472203 496979 472269 496980
rect 470915 496908 470981 496909
rect 470915 496844 470916 496908
rect 470980 496844 470981 496908
rect 470915 496843 470981 496844
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 195244 470414 218898
rect 473514 475174 474134 497940
rect 474414 497181 474474 499530
rect 475702 499530 475828 499590
rect 476040 499590 476100 500106
rect 476992 499590 477052 500106
rect 476040 499530 476130 499590
rect 475702 497725 475762 499530
rect 475699 497724 475765 497725
rect 475699 497660 475700 497724
rect 475764 497660 475765 497724
rect 475699 497659 475765 497660
rect 474411 497180 474477 497181
rect 474411 497116 474412 497180
rect 474476 497116 474477 497180
rect 474411 497115 474477 497116
rect 476070 496909 476130 499530
rect 476990 499530 477052 499590
rect 478080 499590 478140 500106
rect 478488 499590 478548 500106
rect 478080 499530 478154 499590
rect 476990 497725 477050 499530
rect 476987 497724 477053 497725
rect 476987 497660 476988 497724
rect 477052 497660 477053 497724
rect 476987 497659 477053 497660
rect 476067 496908 476133 496909
rect 476067 496844 476068 496908
rect 476132 496844 476133 496908
rect 476067 496843 476133 496844
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 195244 474134 222618
rect 477234 478894 477854 498064
rect 478094 496909 478154 499530
rect 478462 499530 478548 499590
rect 479168 499590 479228 500106
rect 480936 499590 480996 500106
rect 483520 499590 483580 500106
rect 479168 499530 479258 499590
rect 478462 497045 478522 499530
rect 479198 497317 479258 499530
rect 480854 499530 480996 499590
rect 483430 499530 483580 499590
rect 485968 499590 486028 500106
rect 488280 499590 488340 500106
rect 491000 499590 491060 500106
rect 493448 499590 493508 500106
rect 485968 499530 486066 499590
rect 480854 498133 480914 499530
rect 480851 498132 480917 498133
rect 480851 498068 480852 498132
rect 480916 498068 480917 498132
rect 480851 498067 480917 498068
rect 479195 497316 479261 497317
rect 479195 497252 479196 497316
rect 479260 497252 479261 497316
rect 479195 497251 479261 497252
rect 478459 497044 478525 497045
rect 478459 496980 478460 497044
rect 478524 496980 478525 497044
rect 478459 496979 478525 496980
rect 478091 496908 478157 496909
rect 478091 496844 478092 496908
rect 478156 496844 478157 496908
rect 478091 496843 478157 496844
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 195244 477854 226338
rect 480954 482614 481574 497940
rect 483430 496909 483490 499530
rect 483427 496908 483493 496909
rect 483427 496844 483428 496908
rect 483492 496844 483493 496908
rect 483427 496843 483493 496844
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 195244 481574 230058
rect 484674 486334 485294 498064
rect 486006 496909 486066 499530
rect 488214 499530 488340 499590
rect 490974 499530 491060 499590
rect 493366 499530 493508 499590
rect 495896 499590 495956 500106
rect 498480 499590 498540 500106
rect 500928 499590 500988 500106
rect 503512 499590 503572 500106
rect 505960 499590 506020 500106
rect 508544 499590 508604 500106
rect 495896 499530 496002 499590
rect 498480 499530 498578 499590
rect 488214 496909 488274 499530
rect 486003 496908 486069 496909
rect 486003 496844 486004 496908
rect 486068 496844 486069 496908
rect 486003 496843 486069 496844
rect 488211 496908 488277 496909
rect 488211 496844 488212 496908
rect 488276 496844 488277 496908
rect 488211 496843 488277 496844
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484674 450334 485294 485778
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 484674 414334 485294 449778
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 484674 378334 485294 413778
rect 484674 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 485294 378334
rect 484674 378014 485294 378098
rect 484674 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 485294 378014
rect 484674 342334 485294 377778
rect 484674 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 485294 342334
rect 484674 342014 485294 342098
rect 484674 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 485294 342014
rect 484674 306334 485294 341778
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 234334 485294 269778
rect 484674 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 485294 234334
rect 484674 234014 485294 234098
rect 484674 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 485294 234014
rect 484674 198334 485294 233778
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 195244 485294 197778
rect 488394 490054 489014 497940
rect 490974 496909 491034 499530
rect 490971 496908 491037 496909
rect 490971 496844 490972 496908
rect 491036 496844 491037 496908
rect 490971 496843 491037 496844
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454054 489014 489498
rect 488394 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 489014 454054
rect 488394 453734 489014 453818
rect 488394 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 489014 453734
rect 488394 418054 489014 453498
rect 488394 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 489014 418054
rect 488394 417734 489014 417818
rect 488394 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 489014 417734
rect 488394 382054 489014 417498
rect 488394 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 489014 382054
rect 488394 381734 489014 381818
rect 488394 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 489014 381734
rect 488394 346054 489014 381498
rect 488394 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 489014 346054
rect 488394 345734 489014 345818
rect 488394 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 489014 345734
rect 488394 310054 489014 345498
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 238054 489014 273498
rect 488394 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 489014 238054
rect 488394 237734 489014 237818
rect 488394 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 489014 237734
rect 488394 202054 489014 237498
rect 488394 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 489014 202054
rect 488394 201734 489014 201818
rect 488394 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 489014 201734
rect 488394 195244 489014 201498
rect 492114 493774 492734 498064
rect 493366 496909 493426 499530
rect 495942 498133 496002 499530
rect 495939 498132 496005 498133
rect 495939 498068 495940 498132
rect 496004 498068 496005 498132
rect 495939 498067 496005 498068
rect 495834 497494 496454 497940
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 493363 496908 493429 496909
rect 493363 496844 493364 496908
rect 493428 496844 493429 496908
rect 493363 496843 493429 496844
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 492114 385774 492734 421218
rect 492114 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 492734 385774
rect 492114 385454 492734 385538
rect 492114 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 492734 385454
rect 492114 349774 492734 385218
rect 492114 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 492734 349774
rect 492114 349454 492734 349538
rect 492114 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 492734 349454
rect 492114 313774 492734 349218
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 241774 492734 277218
rect 492114 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 492734 241774
rect 492114 241454 492734 241538
rect 492114 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 492734 241454
rect 492114 205774 492734 241218
rect 492114 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 492734 205774
rect 492114 205454 492734 205538
rect 492114 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 492734 205454
rect 492114 195244 492734 205218
rect 495834 461494 496454 496938
rect 498518 496909 498578 499530
rect 500910 499530 500988 499590
rect 503486 499530 503572 499590
rect 505878 499530 506020 499590
rect 508454 499530 508604 499590
rect 510992 499590 511052 500106
rect 513440 499590 513500 500106
rect 515888 499590 515948 500106
rect 518472 499590 518532 500106
rect 510992 499530 511090 499590
rect 500910 496909 500970 499530
rect 503486 496909 503546 499530
rect 505878 498133 505938 499530
rect 505875 498132 505941 498133
rect 505875 498068 505876 498132
rect 505940 498068 505941 498132
rect 505875 498067 505941 498068
rect 498515 496908 498581 496909
rect 498515 496844 498516 496908
rect 498580 496844 498581 496908
rect 498515 496843 498581 496844
rect 500907 496908 500973 496909
rect 500907 496844 500908 496908
rect 500972 496844 500973 496908
rect 500907 496843 500973 496844
rect 503483 496908 503549 496909
rect 503483 496844 503484 496908
rect 503548 496844 503549 496908
rect 503483 496843 503549 496844
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 353494 496454 388938
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 495834 317494 496454 352938
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 245494 496454 280938
rect 495834 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 496454 245494
rect 495834 245174 496454 245258
rect 495834 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 496454 245174
rect 495834 209494 496454 244938
rect 495834 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 496454 209494
rect 495834 209174 496454 209258
rect 495834 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 496454 209174
rect 495834 195244 496454 208938
rect 505794 471454 506414 497940
rect 508454 496909 508514 499530
rect 508451 496908 508517 496909
rect 508451 496844 508452 496908
rect 508516 496844 508517 496908
rect 508451 496843 508517 496844
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 195244 506414 218898
rect 509514 475174 510134 498064
rect 511030 496909 511090 499530
rect 513422 499530 513500 499590
rect 515814 499530 515948 499590
rect 518390 499530 518532 499590
rect 520920 499590 520980 500106
rect 523368 499590 523428 500106
rect 525952 499590 526012 500106
rect 520920 499530 521026 499590
rect 513422 498133 513482 499530
rect 513419 498132 513485 498133
rect 513419 498068 513420 498132
rect 513484 498068 513485 498132
rect 513419 498067 513485 498068
rect 511027 496908 511093 496909
rect 511027 496844 511028 496908
rect 511092 496844 511093 496908
rect 511027 496843 511093 496844
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 195244 510134 222618
rect 513234 478894 513854 497940
rect 515814 496909 515874 499530
rect 515811 496908 515877 496909
rect 515811 496844 515812 496908
rect 515876 496844 515877 496908
rect 515811 496843 515877 496844
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 195244 513854 226338
rect 516954 482614 517574 498064
rect 518390 496909 518450 499530
rect 520966 498133 521026 499530
rect 523358 499530 523428 499590
rect 525934 499530 526012 499590
rect 520963 498132 521029 498133
rect 520963 498068 520964 498132
rect 521028 498068 521029 498132
rect 520963 498067 521029 498068
rect 518387 496908 518453 496909
rect 518387 496844 518388 496908
rect 518452 496844 518453 496908
rect 518387 496843 518453 496844
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 195244 517574 230058
rect 520674 486334 521294 497940
rect 523358 496909 523418 499530
rect 523355 496908 523421 496909
rect 523355 496844 523356 496908
rect 523420 496844 523421 496908
rect 523355 496843 523421 496844
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 234334 521294 269778
rect 520674 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 521294 234334
rect 520674 234014 521294 234098
rect 520674 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 521294 234014
rect 520674 198334 521294 233778
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 195244 521294 197778
rect 524394 490054 525014 498064
rect 525934 496909 525994 499530
rect 525931 496908 525997 496909
rect 525931 496844 525932 496908
rect 525996 496844 525997 496908
rect 525931 496843 525997 496844
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 238054 525014 273498
rect 524394 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 525014 238054
rect 524394 237734 525014 237818
rect 524394 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 525014 237734
rect 524394 202054 525014 237498
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 524394 195244 525014 201498
rect 528114 493774 528734 498064
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 241774 528734 277218
rect 528114 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 528734 241774
rect 528114 241454 528734 241538
rect 528114 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 528734 241454
rect 528114 205774 528734 241218
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 528114 195244 528734 205218
rect 531834 497494 532454 498064
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 531834 195244 532454 208938
rect 541794 471454 542414 498064
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 195244 542414 218898
rect 545514 475174 546134 498064
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 195244 546134 222618
rect 549234 478894 549854 498064
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 195244 549854 226338
rect 552954 482614 553574 498064
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 550955 196076 551021 196077
rect 550955 196012 550956 196076
rect 551020 196012 551021 196076
rect 550955 196011 551021 196012
rect 550958 193490 551018 196011
rect 552954 195244 553574 230058
rect 556674 486334 557294 498064
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 195244 557294 197778
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 550840 193430 551018 193490
rect 550840 193202 550900 193430
rect 420272 187174 420620 187206
rect 420272 186938 420328 187174
rect 420564 186938 420620 187174
rect 420272 186854 420620 186938
rect 420272 186618 420328 186854
rect 420564 186618 420620 186854
rect 420272 186586 420620 186618
rect 556000 187174 556348 187206
rect 556000 186938 556056 187174
rect 556292 186938 556348 187174
rect 556000 186854 556348 186938
rect 556000 186618 556056 186854
rect 556292 186618 556348 186854
rect 556000 186586 556348 186618
rect 420952 183454 421300 183486
rect 420952 183218 421008 183454
rect 421244 183218 421300 183454
rect 420952 183134 421300 183218
rect 420952 182898 421008 183134
rect 421244 182898 421300 183134
rect 420952 182866 421300 182898
rect 555320 183454 555668 183486
rect 555320 183218 555376 183454
rect 555612 183218 555668 183454
rect 555320 183134 555668 183218
rect 555320 182898 555376 183134
rect 555612 182898 555668 183134
rect 555320 182866 555668 182898
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 420272 151174 420620 151206
rect 420272 150938 420328 151174
rect 420564 150938 420620 151174
rect 420272 150854 420620 150938
rect 420272 150618 420328 150854
rect 420564 150618 420620 150854
rect 420272 150586 420620 150618
rect 556000 151174 556348 151206
rect 556000 150938 556056 151174
rect 556292 150938 556348 151174
rect 556000 150854 556348 150938
rect 556000 150618 556056 150854
rect 556292 150618 556348 150854
rect 556000 150586 556348 150618
rect 420952 147454 421300 147486
rect 420952 147218 421008 147454
rect 421244 147218 421300 147454
rect 420952 147134 421300 147218
rect 420952 146898 421008 147134
rect 421244 146898 421300 147134
rect 420952 146866 421300 146898
rect 555320 147454 555668 147486
rect 555320 147218 555376 147454
rect 555612 147218 555668 147454
rect 555320 147134 555668 147218
rect 555320 146898 555376 147134
rect 555612 146898 555668 147134
rect 555320 146866 555668 146898
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 420272 115174 420620 115206
rect 420272 114938 420328 115174
rect 420564 114938 420620 115174
rect 420272 114854 420620 114938
rect 420272 114618 420328 114854
rect 420564 114618 420620 114854
rect 420272 114586 420620 114618
rect 556000 115174 556348 115206
rect 556000 114938 556056 115174
rect 556292 114938 556348 115174
rect 556000 114854 556348 114938
rect 556000 114618 556056 114854
rect 556292 114618 556348 114854
rect 556000 114586 556348 114618
rect 420952 111337 421300 111486
rect 419763 111212 419829 111213
rect 419763 111148 419764 111212
rect 419828 111148 419829 111212
rect 419763 111147 419829 111148
rect 419027 106996 419093 106997
rect 419027 106932 419028 106996
rect 419092 106932 419093 106996
rect 419027 106931 419093 106932
rect 418843 19140 418909 19141
rect 418843 19076 418844 19140
rect 418908 19076 418909 19140
rect 418843 19075 418909 19076
rect 418659 19004 418725 19005
rect 418659 18940 418660 19004
rect 418724 18940 418725 19004
rect 418659 18939 418725 18940
rect 419766 3637 419826 111147
rect 420952 111101 421008 111337
rect 421244 111101 421300 111337
rect 419947 111076 420013 111077
rect 419947 111012 419948 111076
rect 420012 111012 420013 111076
rect 419947 111011 420013 111012
rect 419950 3773 420010 111011
rect 420952 110952 421300 111101
rect 555320 111337 555668 111486
rect 555320 111101 555376 111337
rect 555612 111101 555668 111337
rect 555320 110952 555668 111101
rect 436056 109850 436116 110106
rect 437144 109850 437204 110106
rect 438232 109850 438292 110106
rect 436056 109790 436202 109850
rect 436142 107541 436202 109790
rect 437062 109790 437204 109850
rect 438166 109790 438292 109850
rect 439592 109850 439652 110106
rect 440544 109850 440604 110106
rect 441768 109850 441828 110106
rect 439592 109790 439698 109850
rect 440544 109790 440618 109850
rect 437062 107541 437122 109790
rect 438166 107541 438226 109790
rect 439638 107541 439698 109790
rect 440558 107541 440618 109790
rect 441662 109790 441828 109850
rect 443128 109850 443188 110106
rect 444216 109850 444276 110106
rect 445440 109850 445500 110106
rect 446528 109850 446588 110106
rect 447616 109850 447676 110106
rect 448296 109850 448356 110106
rect 448704 109850 448764 110106
rect 443128 109790 443194 109850
rect 444216 109790 444298 109850
rect 445440 109790 445586 109850
rect 441662 107541 441722 109790
rect 443134 107541 443194 109790
rect 444238 107541 444298 109790
rect 445526 107541 445586 109790
rect 446446 109790 446588 109850
rect 447550 109790 447676 109850
rect 448286 109790 448356 109850
rect 448654 109790 448764 109850
rect 450064 109850 450124 110106
rect 450744 109850 450804 110106
rect 451288 109853 451348 110106
rect 450064 109790 450186 109850
rect 446446 107541 446506 109790
rect 447550 107541 447610 109790
rect 436139 107540 436205 107541
rect 436139 107476 436140 107540
rect 436204 107476 436205 107540
rect 436139 107475 436205 107476
rect 437059 107540 437125 107541
rect 437059 107476 437060 107540
rect 437124 107476 437125 107540
rect 437059 107475 437125 107476
rect 438163 107540 438229 107541
rect 438163 107476 438164 107540
rect 438228 107476 438229 107540
rect 438163 107475 438229 107476
rect 439635 107540 439701 107541
rect 439635 107476 439636 107540
rect 439700 107476 439701 107540
rect 439635 107475 439701 107476
rect 440555 107540 440621 107541
rect 440555 107476 440556 107540
rect 440620 107476 440621 107540
rect 440555 107475 440621 107476
rect 441659 107540 441725 107541
rect 441659 107476 441660 107540
rect 441724 107476 441725 107540
rect 441659 107475 441725 107476
rect 443131 107540 443197 107541
rect 443131 107476 443132 107540
rect 443196 107476 443197 107540
rect 443131 107475 443197 107476
rect 444235 107540 444301 107541
rect 444235 107476 444236 107540
rect 444300 107476 444301 107540
rect 444235 107475 444301 107476
rect 445523 107540 445589 107541
rect 445523 107476 445524 107540
rect 445588 107476 445589 107540
rect 445523 107475 445589 107476
rect 446443 107540 446509 107541
rect 446443 107476 446444 107540
rect 446508 107476 446509 107540
rect 446443 107475 446509 107476
rect 447547 107540 447613 107541
rect 447547 107476 447548 107540
rect 447612 107476 447613 107540
rect 447547 107475 447613 107476
rect 448286 107133 448346 109790
rect 448654 107541 448714 109790
rect 450126 107541 450186 109790
rect 450678 109790 450804 109850
rect 451285 109852 451351 109853
rect 450678 107541 450738 109790
rect 451285 109788 451286 109852
rect 451350 109788 451351 109852
rect 451285 109787 451351 109788
rect 452376 109578 452436 110106
rect 453464 109578 453524 110106
rect 452334 109518 452436 109578
rect 453438 109518 453524 109578
rect 453600 109578 453660 110106
rect 454552 109578 454612 110106
rect 455912 109850 455972 110106
rect 453600 109518 453682 109578
rect 452334 107541 452394 109518
rect 448651 107540 448717 107541
rect 448651 107476 448652 107540
rect 448716 107476 448717 107540
rect 448651 107475 448717 107476
rect 450123 107540 450189 107541
rect 450123 107476 450124 107540
rect 450188 107476 450189 107540
rect 450123 107475 450189 107476
rect 450675 107540 450741 107541
rect 450675 107476 450676 107540
rect 450740 107476 450741 107540
rect 450675 107475 450741 107476
rect 452331 107540 452397 107541
rect 452331 107476 452332 107540
rect 452396 107476 452397 107540
rect 452331 107475 452397 107476
rect 453438 107133 453498 109518
rect 453622 107541 453682 109518
rect 454542 109518 454612 109578
rect 455830 109790 455972 109850
rect 454542 107541 454602 109518
rect 455830 107541 455890 109790
rect 456048 109578 456108 110106
rect 457000 109581 457060 110106
rect 456014 109518 456108 109578
rect 456997 109580 457063 109581
rect 456014 107541 456074 109518
rect 456997 109516 456998 109580
rect 457062 109516 457063 109580
rect 458088 109578 458148 110106
rect 458496 109850 458556 110106
rect 456997 109515 457063 109516
rect 458038 109518 458148 109578
rect 458406 109790 458556 109850
rect 458038 108493 458098 109518
rect 458035 108492 458101 108493
rect 458035 108428 458036 108492
rect 458100 108428 458101 108492
rect 458035 108427 458101 108428
rect 458406 107541 458466 109790
rect 459448 109578 459508 110106
rect 460672 109578 460732 110106
rect 461080 109581 461140 110106
rect 461760 109850 461820 110106
rect 462848 109850 462908 110106
rect 461718 109790 461820 109850
rect 462822 109790 462908 109850
rect 463528 109850 463588 110106
rect 463936 109850 463996 110106
rect 465296 109850 465356 110106
rect 465976 109850 466036 110106
rect 466384 109850 466444 110106
rect 467608 109850 467668 110106
rect 463528 109790 463618 109850
rect 459448 109518 459570 109578
rect 459510 107541 459570 109518
rect 460614 109518 460732 109578
rect 461077 109580 461143 109581
rect 460614 107541 460674 109518
rect 461077 109516 461078 109580
rect 461142 109516 461143 109580
rect 461077 109515 461143 109516
rect 461718 107541 461778 109790
rect 462822 107541 462882 109790
rect 453619 107540 453685 107541
rect 453619 107476 453620 107540
rect 453684 107476 453685 107540
rect 453619 107475 453685 107476
rect 454539 107540 454605 107541
rect 454539 107476 454540 107540
rect 454604 107476 454605 107540
rect 454539 107475 454605 107476
rect 455827 107540 455893 107541
rect 455827 107476 455828 107540
rect 455892 107476 455893 107540
rect 455827 107475 455893 107476
rect 456011 107540 456077 107541
rect 456011 107476 456012 107540
rect 456076 107476 456077 107540
rect 456011 107475 456077 107476
rect 458403 107540 458469 107541
rect 458403 107476 458404 107540
rect 458468 107476 458469 107540
rect 458403 107475 458469 107476
rect 459507 107540 459573 107541
rect 459507 107476 459508 107540
rect 459572 107476 459573 107540
rect 459507 107475 459573 107476
rect 460611 107540 460677 107541
rect 460611 107476 460612 107540
rect 460676 107476 460677 107540
rect 460611 107475 460677 107476
rect 461715 107540 461781 107541
rect 461715 107476 461716 107540
rect 461780 107476 461781 107540
rect 461715 107475 461781 107476
rect 462819 107540 462885 107541
rect 462819 107476 462820 107540
rect 462884 107476 462885 107540
rect 462819 107475 462885 107476
rect 463558 107405 463618 109790
rect 463926 109790 463996 109850
rect 465214 109790 465356 109850
rect 465950 109790 466036 109850
rect 466318 109790 466444 109850
rect 467606 109790 467668 109850
rect 468288 109850 468348 110106
rect 468696 109850 468756 110106
rect 469784 109850 469844 110106
rect 471008 109850 471068 110106
rect 468288 109790 468402 109850
rect 468696 109790 468770 109850
rect 469784 109790 469874 109850
rect 463926 107541 463986 109790
rect 465214 107541 465274 109790
rect 465950 108901 466010 109790
rect 465947 108900 466013 108901
rect 465947 108836 465948 108900
rect 466012 108836 466013 108900
rect 465947 108835 466013 108836
rect 466318 107541 466378 109790
rect 467606 107541 467666 109790
rect 468342 109173 468402 109790
rect 468339 109172 468405 109173
rect 468339 109108 468340 109172
rect 468404 109108 468405 109172
rect 468339 109107 468405 109108
rect 468710 107541 468770 109790
rect 469814 107541 469874 109790
rect 470918 109790 471068 109850
rect 471144 109850 471204 110106
rect 472232 109850 472292 110106
rect 473320 109850 473380 110106
rect 473592 109850 473652 110106
rect 471144 109790 471346 109850
rect 470918 109037 470978 109790
rect 470915 109036 470981 109037
rect 470915 108972 470916 109036
rect 470980 108972 470981 109036
rect 470915 108971 470981 108972
rect 471286 107541 471346 109790
rect 472206 109790 472292 109850
rect 473310 109790 473380 109850
rect 473494 109790 473652 109850
rect 474408 109850 474468 110106
rect 475768 109850 475828 110106
rect 474408 109790 474474 109850
rect 472206 107541 472266 109790
rect 473310 107541 473370 109790
rect 463923 107540 463989 107541
rect 463923 107476 463924 107540
rect 463988 107476 463989 107540
rect 463923 107475 463989 107476
rect 465211 107540 465277 107541
rect 465211 107476 465212 107540
rect 465276 107476 465277 107540
rect 465211 107475 465277 107476
rect 466315 107540 466381 107541
rect 466315 107476 466316 107540
rect 466380 107476 466381 107540
rect 466315 107475 466381 107476
rect 467603 107540 467669 107541
rect 467603 107476 467604 107540
rect 467668 107476 467669 107540
rect 467603 107475 467669 107476
rect 468707 107540 468773 107541
rect 468707 107476 468708 107540
rect 468772 107476 468773 107540
rect 468707 107475 468773 107476
rect 469811 107540 469877 107541
rect 469811 107476 469812 107540
rect 469876 107476 469877 107540
rect 469811 107475 469877 107476
rect 471283 107540 471349 107541
rect 471283 107476 471284 107540
rect 471348 107476 471349 107540
rect 471283 107475 471349 107476
rect 472203 107540 472269 107541
rect 472203 107476 472204 107540
rect 472268 107476 472269 107540
rect 472203 107475 472269 107476
rect 473307 107540 473373 107541
rect 473307 107476 473308 107540
rect 473372 107476 473373 107540
rect 473307 107475 473373 107476
rect 463555 107404 463621 107405
rect 463555 107340 463556 107404
rect 463620 107340 463621 107404
rect 463555 107339 463621 107340
rect 448283 107132 448349 107133
rect 448283 107068 448284 107132
rect 448348 107068 448349 107132
rect 448283 107067 448349 107068
rect 453435 107132 453501 107133
rect 453435 107068 453436 107132
rect 453500 107068 453501 107132
rect 453435 107067 453501 107068
rect 473494 106997 473554 109790
rect 474414 107541 474474 109790
rect 475702 109790 475828 109850
rect 476040 109850 476100 110106
rect 476992 109850 477052 110106
rect 476040 109790 476130 109850
rect 475702 107541 475762 109790
rect 476070 109717 476130 109790
rect 476990 109790 477052 109850
rect 478080 109850 478140 110106
rect 478488 109850 478548 110106
rect 478080 109790 478154 109850
rect 476067 109716 476133 109717
rect 476067 109652 476068 109716
rect 476132 109652 476133 109716
rect 476067 109651 476133 109652
rect 474411 107540 474477 107541
rect 474411 107476 474412 107540
rect 474476 107476 474477 107540
rect 474411 107475 474477 107476
rect 475699 107540 475765 107541
rect 475699 107476 475700 107540
rect 475764 107476 475765 107540
rect 475699 107475 475765 107476
rect 476990 107133 477050 109790
rect 478094 107541 478154 109790
rect 478462 109790 478548 109850
rect 479168 109850 479228 110106
rect 480936 109853 480996 110106
rect 483520 109853 483580 110106
rect 485968 109853 486028 110106
rect 488280 109853 488340 110106
rect 491000 109853 491060 110106
rect 480933 109852 480999 109853
rect 479168 109790 479258 109850
rect 478091 107540 478157 107541
rect 478091 107476 478092 107540
rect 478156 107476 478157 107540
rect 478091 107475 478157 107476
rect 478462 107269 478522 109790
rect 479198 107541 479258 109790
rect 480933 109788 480934 109852
rect 480998 109788 480999 109852
rect 480933 109787 480999 109788
rect 483517 109852 483583 109853
rect 483517 109788 483518 109852
rect 483582 109788 483583 109852
rect 483517 109787 483583 109788
rect 485965 109852 486031 109853
rect 485965 109788 485966 109852
rect 486030 109788 486031 109852
rect 485965 109787 486031 109788
rect 488277 109852 488343 109853
rect 488277 109788 488278 109852
rect 488342 109788 488343 109852
rect 488277 109787 488343 109788
rect 490997 109852 491063 109853
rect 490997 109788 490998 109852
rect 491062 109788 491063 109852
rect 490997 109787 491063 109788
rect 493448 109717 493508 110106
rect 495896 109717 495956 110106
rect 498480 109717 498540 110106
rect 500928 109850 500988 110106
rect 503512 109850 503572 110106
rect 500910 109790 500988 109850
rect 503486 109790 503572 109850
rect 493445 109716 493511 109717
rect 493445 109652 493446 109716
rect 493510 109652 493511 109716
rect 493445 109651 493511 109652
rect 495893 109716 495959 109717
rect 495893 109652 495894 109716
rect 495958 109652 495959 109716
rect 495893 109651 495959 109652
rect 498477 109716 498543 109717
rect 498477 109652 498478 109716
rect 498542 109652 498543 109716
rect 498477 109651 498543 109652
rect 500910 109037 500970 109790
rect 503486 109037 503546 109790
rect 505960 109581 506020 110106
rect 508544 109581 508604 110106
rect 510992 109850 511052 110106
rect 513440 109850 513500 110106
rect 510992 109790 511090 109850
rect 505957 109580 506023 109581
rect 505957 109516 505958 109580
rect 506022 109516 506023 109580
rect 505957 109515 506023 109516
rect 508541 109580 508607 109581
rect 508541 109516 508542 109580
rect 508606 109516 508607 109580
rect 508541 109515 508607 109516
rect 500907 109036 500973 109037
rect 500907 108972 500908 109036
rect 500972 108972 500973 109036
rect 500907 108971 500973 108972
rect 503483 109036 503549 109037
rect 503483 108972 503484 109036
rect 503548 108972 503549 109036
rect 503483 108971 503549 108972
rect 479195 107540 479261 107541
rect 479195 107476 479196 107540
rect 479260 107476 479261 107540
rect 479195 107475 479261 107476
rect 478459 107268 478525 107269
rect 478459 107204 478460 107268
rect 478524 107204 478525 107268
rect 478459 107203 478525 107204
rect 476987 107132 477053 107133
rect 476987 107068 476988 107132
rect 477052 107068 477053 107132
rect 476987 107067 477053 107068
rect 473491 106996 473557 106997
rect 473491 106932 473492 106996
rect 473556 106932 473557 106996
rect 473491 106931 473557 106932
rect 511030 106725 511090 109790
rect 513422 109790 513500 109850
rect 513422 109037 513482 109790
rect 515888 109581 515948 110106
rect 518472 109581 518532 110106
rect 520920 109850 520980 110106
rect 523368 109850 523428 110106
rect 525952 109850 526012 110106
rect 520920 109790 521026 109850
rect 515885 109580 515951 109581
rect 515885 109516 515886 109580
rect 515950 109516 515951 109580
rect 515885 109515 515951 109516
rect 518469 109580 518535 109581
rect 518469 109516 518470 109580
rect 518534 109516 518535 109580
rect 518469 109515 518535 109516
rect 520966 109037 521026 109790
rect 523358 109790 523428 109850
rect 525934 109790 526012 109850
rect 523358 109037 523418 109790
rect 525934 109037 525994 109790
rect 513419 109036 513485 109037
rect 513419 108972 513420 109036
rect 513484 108972 513485 109036
rect 513419 108971 513485 108972
rect 520963 109036 521029 109037
rect 520963 108972 520964 109036
rect 521028 108972 521029 109036
rect 520963 108971 521029 108972
rect 523355 109036 523421 109037
rect 523355 108972 523356 109036
rect 523420 108972 523421 109036
rect 523355 108971 523421 108972
rect 525931 109036 525997 109037
rect 525931 108972 525932 109036
rect 525996 108972 525997 109036
rect 525931 108971 525997 108972
rect 511027 106724 511093 106725
rect 511027 106660 511028 106724
rect 511092 106660 511093 106724
rect 511027 106659 511093 106660
rect 550771 105364 550837 105365
rect 550771 105300 550772 105364
rect 550836 105300 550837 105364
rect 550771 105299 550837 105300
rect 550774 103530 550834 105299
rect 550774 103470 550900 103530
rect 550840 103202 550900 103470
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 420272 79174 420620 79206
rect 420272 78938 420328 79174
rect 420564 78938 420620 79174
rect 420272 78854 420620 78938
rect 420272 78618 420328 78854
rect 420564 78618 420620 78854
rect 420272 78586 420620 78618
rect 556000 79174 556348 79206
rect 556000 78938 556056 79174
rect 556292 78938 556348 79174
rect 556000 78854 556348 78938
rect 556000 78618 556056 78854
rect 556292 78618 556348 78854
rect 556000 78586 556348 78618
rect 420952 75454 421300 75486
rect 420952 75218 421008 75454
rect 421244 75218 421300 75454
rect 420952 75134 421300 75218
rect 420952 74898 421008 75134
rect 421244 74898 421300 75134
rect 420952 74866 421300 74898
rect 555320 75454 555668 75486
rect 555320 75218 555376 75454
rect 555612 75218 555668 75454
rect 555320 75134 555668 75218
rect 555320 74898 555376 75134
rect 555612 74898 555668 75134
rect 555320 74866 555668 74898
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 420272 43174 420620 43206
rect 420272 42938 420328 43174
rect 420564 42938 420620 43174
rect 420272 42854 420620 42938
rect 420272 42618 420328 42854
rect 420564 42618 420620 42854
rect 420272 42586 420620 42618
rect 556000 43174 556348 43206
rect 556000 42938 556056 43174
rect 556292 42938 556348 43174
rect 556000 42854 556348 42938
rect 556000 42618 556056 42854
rect 556292 42618 556348 42854
rect 556000 42586 556348 42618
rect 420952 39454 421300 39486
rect 420952 39218 421008 39454
rect 421244 39218 421300 39454
rect 420952 39134 421300 39218
rect 420952 38898 421008 39134
rect 421244 38898 421300 39134
rect 420952 38866 421300 38898
rect 555320 39454 555668 39486
rect 555320 39218 555376 39454
rect 555612 39218 555668 39454
rect 555320 39134 555668 39218
rect 555320 38898 555376 39134
rect 555612 38898 555668 39134
rect 555320 38866 555668 38898
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 436056 19410 436116 20060
rect 437144 19410 437204 20060
rect 436056 19350 436202 19410
rect 419947 3772 420013 3773
rect 419947 3708 419948 3772
rect 420012 3708 420013 3772
rect 419947 3707 420013 3708
rect 419763 3636 419829 3637
rect 419763 3572 419764 3636
rect 419828 3572 419829 3636
rect 419763 3571 419829 3572
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 433794 3454 434414 18064
rect 436142 17917 436202 19350
rect 437062 19350 437204 19410
rect 438232 19410 438292 20060
rect 439592 19410 439652 20060
rect 440544 19410 440604 20060
rect 441768 19410 441828 20060
rect 443128 19410 443188 20060
rect 444216 19410 444276 20060
rect 445440 19410 445500 20060
rect 446528 19410 446588 20060
rect 447616 19685 447676 20060
rect 447613 19684 447679 19685
rect 447613 19620 447614 19684
rect 447678 19620 447679 19684
rect 447613 19619 447679 19620
rect 448296 19410 448356 20060
rect 448704 19685 448764 20060
rect 450064 19685 450124 20060
rect 448701 19684 448767 19685
rect 448701 19620 448702 19684
rect 448766 19620 448767 19684
rect 448701 19619 448767 19620
rect 450061 19684 450127 19685
rect 450061 19620 450062 19684
rect 450126 19620 450127 19684
rect 450061 19619 450127 19620
rect 450744 19410 450804 20060
rect 451288 19546 451348 20060
rect 452376 19546 452436 20060
rect 453464 19546 453524 20060
rect 451288 19486 451474 19546
rect 438232 19350 438410 19410
rect 439592 19350 439698 19410
rect 440544 19350 440618 19410
rect 441768 19350 442090 19410
rect 443128 19350 443194 19410
rect 444216 19350 444298 19410
rect 445440 19350 445770 19410
rect 437062 17917 437122 19350
rect 436139 17916 436205 17917
rect 436139 17852 436140 17916
rect 436204 17852 436205 17916
rect 436139 17851 436205 17852
rect 437059 17916 437125 17917
rect 437059 17852 437060 17916
rect 437124 17852 437125 17916
rect 437059 17851 437125 17852
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 18064
rect 438350 17917 438410 19350
rect 439638 17917 439698 19350
rect 440558 17917 440618 19350
rect 438347 17916 438413 17917
rect 438347 17852 438348 17916
rect 438412 17852 438413 17916
rect 438347 17851 438413 17852
rect 439635 17916 439701 17917
rect 439635 17852 439636 17916
rect 439700 17852 439701 17916
rect 439635 17851 439701 17852
rect 440555 17916 440621 17917
rect 440555 17852 440556 17916
rect 440620 17852 440621 17916
rect 440555 17851 440621 17852
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 17940
rect 442030 17917 442090 19350
rect 443134 17917 443194 19350
rect 444238 17917 444298 19350
rect 442027 17916 442093 17917
rect 442027 17852 442028 17916
rect 442092 17852 442093 17916
rect 442027 17851 442093 17852
rect 443131 17916 443197 17917
rect 443131 17852 443132 17916
rect 443196 17852 443197 17916
rect 443131 17851 443197 17852
rect 444235 17916 444301 17917
rect 444235 17852 444236 17916
rect 444300 17852 444301 17916
rect 444235 17851 444301 17852
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 14614 445574 17940
rect 445710 17917 445770 19350
rect 446446 19350 446588 19410
rect 448286 19350 448356 19410
rect 450678 19350 450804 19410
rect 446446 17917 446506 19350
rect 448286 17917 448346 19350
rect 445707 17916 445773 17917
rect 445707 17852 445708 17916
rect 445772 17852 445773 17916
rect 445707 17851 445773 17852
rect 446443 17916 446509 17917
rect 446443 17852 446444 17916
rect 446508 17852 446509 17916
rect 446443 17851 446509 17852
rect 448283 17916 448349 17917
rect 448283 17852 448284 17916
rect 448348 17852 448349 17916
rect 448283 17851 448349 17852
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 -4186 449294 17940
rect 450678 17917 450738 19350
rect 451414 17917 451474 19486
rect 452334 19486 452436 19546
rect 453438 19486 453524 19546
rect 453600 19546 453660 20060
rect 454552 19546 454612 20060
rect 455912 19685 455972 20060
rect 455909 19684 455975 19685
rect 455909 19620 455910 19684
rect 455974 19620 455975 19684
rect 455909 19619 455975 19620
rect 456048 19546 456108 20060
rect 453600 19486 453682 19546
rect 452334 17917 452394 19486
rect 453438 17917 453498 19486
rect 450675 17916 450741 17917
rect 450675 17852 450676 17916
rect 450740 17852 450741 17916
rect 450675 17851 450741 17852
rect 451411 17916 451477 17917
rect 451411 17852 451412 17916
rect 451476 17852 451477 17916
rect 451411 17851 451477 17852
rect 452331 17916 452397 17917
rect 452331 17852 452332 17916
rect 452396 17852 452397 17916
rect 452331 17851 452397 17852
rect 453435 17916 453501 17917
rect 453435 17852 453436 17916
rect 453500 17852 453501 17916
rect 453435 17851 453501 17852
rect 453622 16965 453682 19486
rect 454542 19486 454612 19546
rect 456014 19486 456108 19546
rect 457000 19546 457060 20060
rect 458088 19546 458148 20060
rect 458496 19546 458556 20060
rect 459448 19546 459508 20060
rect 460672 19821 460732 20060
rect 460669 19820 460735 19821
rect 460669 19756 460670 19820
rect 460734 19756 460735 19820
rect 460669 19755 460735 19756
rect 461080 19549 461140 20060
rect 461760 19682 461820 20060
rect 462848 19682 462908 20060
rect 461718 19622 461820 19682
rect 462822 19622 462908 19682
rect 463528 19682 463588 20060
rect 463936 19682 463996 20060
rect 465296 19682 465356 20060
rect 465976 19682 466036 20060
rect 466384 19682 466444 20060
rect 467608 19682 467668 20060
rect 463528 19622 463618 19682
rect 457000 19486 457178 19546
rect 454542 17917 454602 19486
rect 456014 17917 456074 19486
rect 457118 17917 457178 19486
rect 458038 19486 458148 19546
rect 458406 19486 458556 19546
rect 459326 19486 459508 19546
rect 461077 19548 461143 19549
rect 458038 17917 458098 19486
rect 458406 18053 458466 19486
rect 458403 18052 458469 18053
rect 458403 17988 458404 18052
rect 458468 17988 458469 18052
rect 458403 17987 458469 17988
rect 459326 17917 459386 19486
rect 461077 19484 461078 19548
rect 461142 19484 461143 19548
rect 461077 19483 461143 19484
rect 461718 17917 461778 19622
rect 462822 17917 462882 19622
rect 463558 18597 463618 19622
rect 463926 19622 463996 19682
rect 465214 19622 465356 19682
rect 465950 19622 466036 19682
rect 466318 19622 466444 19682
rect 467606 19622 467668 19682
rect 463555 18596 463621 18597
rect 463555 18532 463556 18596
rect 463620 18532 463621 18596
rect 463555 18531 463621 18532
rect 463926 17917 463986 19622
rect 454539 17916 454605 17917
rect 454539 17852 454540 17916
rect 454604 17852 454605 17916
rect 454539 17851 454605 17852
rect 456011 17916 456077 17917
rect 456011 17852 456012 17916
rect 456076 17852 456077 17916
rect 456011 17851 456077 17852
rect 457115 17916 457181 17917
rect 457115 17852 457116 17916
rect 457180 17852 457181 17916
rect 457115 17851 457181 17852
rect 458035 17916 458101 17917
rect 458035 17852 458036 17916
rect 458100 17852 458101 17916
rect 458035 17851 458101 17852
rect 459323 17916 459389 17917
rect 459323 17852 459324 17916
rect 459388 17852 459389 17916
rect 459323 17851 459389 17852
rect 461715 17916 461781 17917
rect 461715 17852 461716 17916
rect 461780 17852 461781 17916
rect 461715 17851 461781 17852
rect 462819 17916 462885 17917
rect 462819 17852 462820 17916
rect 462884 17852 462885 17916
rect 462819 17851 462885 17852
rect 463923 17916 463989 17917
rect 463923 17852 463924 17916
rect 463988 17852 463989 17916
rect 463923 17851 463989 17852
rect 465214 17101 465274 19622
rect 465950 18869 466010 19622
rect 465947 18868 466013 18869
rect 465947 18804 465948 18868
rect 466012 18804 466013 18868
rect 465947 18803 466013 18804
rect 466318 17917 466378 19622
rect 467606 17917 467666 19622
rect 468288 19549 468348 20060
rect 468696 19682 468756 20060
rect 469784 19682 469844 20060
rect 468696 19622 468770 19682
rect 468285 19548 468351 19549
rect 468285 19484 468286 19548
rect 468350 19484 468351 19548
rect 468285 19483 468351 19484
rect 468710 17917 468770 19622
rect 469630 19622 469844 19682
rect 466315 17916 466381 17917
rect 466315 17852 466316 17916
rect 466380 17852 466381 17916
rect 466315 17851 466381 17852
rect 467603 17916 467669 17917
rect 467603 17852 467604 17916
rect 467668 17852 467669 17916
rect 467603 17851 467669 17852
rect 468707 17916 468773 17917
rect 468707 17852 468708 17916
rect 468772 17852 468773 17916
rect 468707 17851 468773 17852
rect 469630 17101 469690 19622
rect 471008 19410 471068 20060
rect 470918 19350 471068 19410
rect 471144 19410 471204 20060
rect 472232 19410 472292 20060
rect 473320 19685 473380 20060
rect 473317 19684 473383 19685
rect 473317 19620 473318 19684
rect 473382 19620 473383 19684
rect 473317 19619 473383 19620
rect 473592 19410 473652 20060
rect 471144 19350 471346 19410
rect 470918 18869 470978 19350
rect 470915 18868 470981 18869
rect 470915 18804 470916 18868
rect 470980 18804 470981 18868
rect 470915 18803 470981 18804
rect 465211 17100 465277 17101
rect 465211 17036 465212 17100
rect 465276 17036 465277 17100
rect 465211 17035 465277 17036
rect 469627 17100 469693 17101
rect 469627 17036 469628 17100
rect 469692 17036 469693 17100
rect 469627 17035 469693 17036
rect 453619 16964 453685 16965
rect 453619 16900 453620 16964
rect 453684 16900 453685 16964
rect 453619 16899 453685 16900
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 469794 3454 470414 17940
rect 471286 16829 471346 19350
rect 472206 19350 472292 19410
rect 473310 19350 473652 19410
rect 474408 19410 474468 20060
rect 475768 19410 475828 20060
rect 474408 19350 474474 19410
rect 472206 17237 472266 19350
rect 473310 17781 473370 19350
rect 473307 17780 473373 17781
rect 473307 17716 473308 17780
rect 473372 17716 473373 17780
rect 473307 17715 473373 17716
rect 472203 17236 472269 17237
rect 472203 17172 472204 17236
rect 472268 17172 472269 17236
rect 472203 17171 472269 17172
rect 471283 16828 471349 16829
rect 471283 16764 471284 16828
rect 471348 16764 471349 16828
rect 471283 16763 471349 16764
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 7174 474134 17940
rect 474414 17917 474474 19350
rect 475702 19350 475828 19410
rect 476040 19410 476100 20060
rect 476992 19410 477052 20060
rect 476040 19350 476130 19410
rect 474411 17916 474477 17917
rect 474411 17852 474412 17916
rect 474476 17852 474477 17916
rect 474411 17851 474477 17852
rect 475702 17237 475762 19350
rect 476070 17373 476130 19350
rect 476990 19350 477052 19410
rect 478080 19410 478140 20060
rect 478488 19410 478548 20060
rect 478080 19350 478154 19410
rect 476990 17917 477050 19350
rect 476987 17916 477053 17917
rect 476987 17852 476988 17916
rect 477052 17852 477053 17916
rect 476987 17851 477053 17852
rect 476067 17372 476133 17373
rect 476067 17308 476068 17372
rect 476132 17308 476133 17372
rect 476067 17307 476133 17308
rect 475699 17236 475765 17237
rect 475699 17172 475700 17236
rect 475764 17172 475765 17236
rect 475699 17171 475765 17172
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 10894 477854 18064
rect 478094 16965 478154 19350
rect 478462 19350 478548 19410
rect 479168 19410 479228 20060
rect 480936 19410 480996 20060
rect 483520 19410 483580 20060
rect 485968 19549 486028 20060
rect 488280 19821 488340 20060
rect 488277 19820 488343 19821
rect 488277 19756 488278 19820
rect 488342 19756 488343 19820
rect 488277 19755 488343 19756
rect 491000 19685 491060 20060
rect 493448 19685 493508 20060
rect 490997 19684 491063 19685
rect 490997 19620 490998 19684
rect 491062 19620 491063 19684
rect 490997 19619 491063 19620
rect 493445 19684 493511 19685
rect 493445 19620 493446 19684
rect 493510 19620 493511 19684
rect 493445 19619 493511 19620
rect 495896 19549 495956 20060
rect 485965 19548 486031 19549
rect 485965 19484 485966 19548
rect 486030 19484 486031 19548
rect 485965 19483 486031 19484
rect 495893 19548 495959 19549
rect 495893 19484 495894 19548
rect 495958 19484 495959 19548
rect 495893 19483 495959 19484
rect 479168 19350 479258 19410
rect 478462 17101 478522 19350
rect 479198 17917 479258 19350
rect 480670 19350 480996 19410
rect 483430 19350 483580 19410
rect 498480 19410 498540 20060
rect 500928 19549 500988 20060
rect 503512 19549 503572 20060
rect 500925 19548 500991 19549
rect 500925 19484 500926 19548
rect 500990 19484 500991 19548
rect 500925 19483 500991 19484
rect 503509 19548 503575 19549
rect 503509 19484 503510 19548
rect 503574 19484 503575 19548
rect 503509 19483 503575 19484
rect 505960 19410 506020 20060
rect 508544 19410 508604 20060
rect 498480 19350 498578 19410
rect 479195 17916 479261 17917
rect 479195 17852 479196 17916
rect 479260 17852 479261 17916
rect 479195 17851 479261 17852
rect 480670 17781 480730 19350
rect 480667 17780 480733 17781
rect 480667 17716 480668 17780
rect 480732 17716 480733 17780
rect 480667 17715 480733 17716
rect 478459 17100 478525 17101
rect 478459 17036 478460 17100
rect 478524 17036 478525 17100
rect 478459 17035 478525 17036
rect 478091 16964 478157 16965
rect 478091 16900 478092 16964
rect 478156 16900 478157 16964
rect 478091 16899 478157 16900
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 14614 481574 17940
rect 483430 17645 483490 19350
rect 498518 19277 498578 19350
rect 505878 19350 506020 19410
rect 508454 19350 508604 19410
rect 510992 19410 511052 20060
rect 513440 19410 513500 20060
rect 515888 19410 515948 20060
rect 518472 19410 518532 20060
rect 510992 19350 511090 19410
rect 498515 19276 498581 19277
rect 498515 19212 498516 19276
rect 498580 19212 498581 19276
rect 498515 19211 498581 19212
rect 505878 18869 505938 19350
rect 508454 18869 508514 19350
rect 505875 18868 505941 18869
rect 505875 18804 505876 18868
rect 505940 18804 505941 18868
rect 505875 18803 505941 18804
rect 508451 18868 508517 18869
rect 508451 18804 508452 18868
rect 508516 18804 508517 18868
rect 508451 18803 508517 18804
rect 484674 18023 485294 18064
rect 484674 17787 484706 18023
rect 484942 17787 485026 18023
rect 485262 17787 485294 18023
rect 483427 17644 483493 17645
rect 483427 17580 483428 17644
rect 483492 17580 483493 17644
rect 483427 17579 483493 17580
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 -4186 485294 17787
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 505794 3454 506414 17940
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 7174 510134 18064
rect 511030 16693 511090 19350
rect 513422 19350 513500 19410
rect 515814 19350 515948 19410
rect 518390 19350 518532 19410
rect 520920 19410 520980 20060
rect 523368 19410 523428 20060
rect 525952 19410 526012 20060
rect 520920 19350 521026 19410
rect 513422 19005 513482 19350
rect 515814 19005 515874 19350
rect 518390 19141 518450 19350
rect 520966 19277 521026 19350
rect 523358 19350 523428 19410
rect 525934 19350 526012 19410
rect 520963 19276 521029 19277
rect 520963 19212 520964 19276
rect 521028 19212 521029 19276
rect 520963 19211 521029 19212
rect 518387 19140 518453 19141
rect 518387 19076 518388 19140
rect 518452 19076 518453 19140
rect 518387 19075 518453 19076
rect 513419 19004 513485 19005
rect 513419 18940 513420 19004
rect 513484 18940 513485 19004
rect 513419 18939 513485 18940
rect 515811 19004 515877 19005
rect 515811 18940 515812 19004
rect 515876 18940 515877 19004
rect 515811 18939 515877 18940
rect 523358 18733 523418 19350
rect 525934 18733 525994 19350
rect 523355 18732 523421 18733
rect 523355 18668 523356 18732
rect 523420 18668 523421 18732
rect 523355 18667 523421 18668
rect 525931 18732 525997 18733
rect 525931 18668 525932 18732
rect 525996 18668 525997 18732
rect 525931 18667 525997 18668
rect 511027 16692 511093 16693
rect 511027 16628 511028 16692
rect 511092 16628 511093 16692
rect 511027 16627 511093 16628
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 10894 513854 17940
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 14614 517574 18064
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 -4186 521294 17940
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 541794 3454 542414 18064
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 18064
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 18064
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 18064
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18023 557294 18064
rect 556674 17787 556706 18023
rect 556942 17787 557026 18023
rect 557262 17787 557294 18023
rect 556674 -4186 557294 17787
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 20328 654938 20564 655174
rect 20328 654618 20564 654854
rect 156056 654938 156292 655174
rect 156056 654618 156292 654854
rect 21008 651218 21244 651454
rect 21008 650898 21244 651134
rect 155376 651218 155612 651454
rect 155376 650898 155612 651134
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 20328 618938 20564 619174
rect 20328 618618 20564 618854
rect 156056 618938 156292 619174
rect 156056 618618 156292 618854
rect 21008 615218 21244 615454
rect 21008 614898 21244 615134
rect 155376 615218 155612 615454
rect 155376 614898 155612 615134
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 160706 594098 160942 594334
rect 161026 594098 161262 594334
rect 160706 593778 160942 594014
rect 161026 593778 161262 594014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 20328 582693 20564 582929
rect 156056 582693 156292 582929
rect 21008 579218 21244 579454
rect 21008 578898 21244 579134
rect 155376 579218 155612 579454
rect 155376 578898 155612 579134
rect 160706 558098 160942 558334
rect 161026 558098 161262 558334
rect 160706 557778 160942 558014
rect 161026 557778 161262 558014
rect 20328 546938 20564 547174
rect 20328 546618 20564 546854
rect 156056 546938 156292 547174
rect 156056 546618 156292 546854
rect 21008 543218 21244 543454
rect 21008 542898 21244 543134
rect 155376 543218 155612 543454
rect 155376 542898 155612 543134
rect 160706 522098 160942 522334
rect 161026 522098 161262 522334
rect 160706 521778 160942 522014
rect 161026 521778 161262 522014
rect 20328 510938 20564 511174
rect 20328 510618 20564 510854
rect 156056 510938 156292 511174
rect 156056 510618 156292 510854
rect 21008 507218 21244 507454
rect 21008 506898 21244 507134
rect 155376 507218 155612 507454
rect 155376 506898 155612 507134
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 63866 497258 64102 497494
rect 64186 497258 64422 497494
rect 63866 496938 64102 497174
rect 64186 496938 64422 497174
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 60146 241538 60382 241774
rect 60466 241538 60702 241774
rect 60146 241218 60382 241454
rect 60466 241218 60702 241454
rect 60146 205538 60382 205774
rect 60466 205538 60702 205774
rect 60146 205218 60382 205454
rect 60466 205218 60702 205454
rect 63866 461258 64102 461494
rect 64186 461258 64422 461494
rect 63866 460938 64102 461174
rect 64186 460938 64422 461174
rect 63866 425258 64102 425494
rect 64186 425258 64422 425494
rect 63866 424938 64102 425174
rect 64186 424938 64422 425174
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 63866 317258 64102 317494
rect 64186 317258 64422 317494
rect 63866 316938 64102 317174
rect 64186 316938 64422 317174
rect 63866 281258 64102 281494
rect 64186 281258 64422 281494
rect 63866 280938 64102 281174
rect 64186 280938 64422 281174
rect 63866 245258 64102 245494
rect 64186 245258 64422 245494
rect 63866 244938 64102 245174
rect 64186 244938 64422 245174
rect 63866 209258 64102 209494
rect 64186 209258 64422 209494
rect 63866 208938 64102 209174
rect 64186 208938 64422 209174
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 88706 486098 88942 486334
rect 89026 486098 89262 486334
rect 88706 485778 88942 486014
rect 89026 485778 89262 486014
rect 88706 450098 88942 450334
rect 89026 450098 89262 450334
rect 88706 449778 88942 450014
rect 89026 449778 89262 450014
rect 88706 414098 88942 414334
rect 89026 414098 89262 414334
rect 88706 413778 88942 414014
rect 89026 413778 89262 414014
rect 88706 378098 88942 378334
rect 89026 378098 89262 378334
rect 88706 377778 88942 378014
rect 89026 377778 89262 378014
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 88706 306098 88942 306334
rect 89026 306098 89262 306334
rect 88706 305778 88942 306014
rect 89026 305778 89262 306014
rect 88706 270098 88942 270334
rect 89026 270098 89262 270334
rect 88706 269778 88942 270014
rect 89026 269778 89262 270014
rect 88706 234098 88942 234334
rect 89026 234098 89262 234334
rect 88706 233778 88942 234014
rect 89026 233778 89262 234014
rect 88706 198098 88942 198334
rect 89026 198098 89262 198334
rect 88706 197778 88942 198014
rect 89026 197778 89262 198014
rect 92426 489818 92662 490054
rect 92746 489818 92982 490054
rect 92426 489498 92662 489734
rect 92746 489498 92982 489734
rect 92426 453818 92662 454054
rect 92746 453818 92982 454054
rect 92426 453498 92662 453734
rect 92746 453498 92982 453734
rect 92426 417818 92662 418054
rect 92746 417818 92982 418054
rect 92426 417498 92662 417734
rect 92746 417498 92982 417734
rect 92426 381818 92662 382054
rect 92746 381818 92982 382054
rect 92426 381498 92662 381734
rect 92746 381498 92982 381734
rect 92426 345818 92662 346054
rect 92746 345818 92982 346054
rect 92426 345498 92662 345734
rect 92746 345498 92982 345734
rect 92426 309818 92662 310054
rect 92746 309818 92982 310054
rect 92426 309498 92662 309734
rect 92746 309498 92982 309734
rect 92426 273818 92662 274054
rect 92746 273818 92982 274054
rect 92426 273498 92662 273734
rect 92746 273498 92982 273734
rect 92426 237818 92662 238054
rect 92746 237818 92982 238054
rect 92426 237498 92662 237734
rect 92746 237498 92982 237734
rect 92426 201818 92662 202054
rect 92746 201818 92982 202054
rect 92426 201498 92662 201734
rect 92746 201498 92982 201734
rect 99866 497258 100102 497494
rect 100186 497258 100422 497494
rect 99866 496938 100102 497174
rect 100186 496938 100422 497174
rect 96146 493538 96382 493774
rect 96466 493538 96702 493774
rect 96146 493218 96382 493454
rect 96466 493218 96702 493454
rect 96146 457538 96382 457774
rect 96466 457538 96702 457774
rect 96146 457218 96382 457454
rect 96466 457218 96702 457454
rect 96146 421538 96382 421774
rect 96466 421538 96702 421774
rect 96146 421218 96382 421454
rect 96466 421218 96702 421454
rect 96146 385538 96382 385774
rect 96466 385538 96702 385774
rect 96146 385218 96382 385454
rect 96466 385218 96702 385454
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 96146 313538 96382 313774
rect 96466 313538 96702 313774
rect 96146 313218 96382 313454
rect 96466 313218 96702 313454
rect 96146 277538 96382 277774
rect 96466 277538 96702 277774
rect 96146 277218 96382 277454
rect 96466 277218 96702 277454
rect 96146 241538 96382 241774
rect 96466 241538 96702 241774
rect 96146 241218 96382 241454
rect 96466 241218 96702 241454
rect 96146 205538 96382 205774
rect 96466 205538 96702 205774
rect 96146 205218 96382 205454
rect 96466 205218 96702 205454
rect 99866 461258 100102 461494
rect 100186 461258 100422 461494
rect 99866 460938 100102 461174
rect 100186 460938 100422 461174
rect 99866 425258 100102 425494
rect 100186 425258 100422 425494
rect 99866 424938 100102 425174
rect 100186 424938 100422 425174
rect 99866 389258 100102 389494
rect 100186 389258 100422 389494
rect 99866 388938 100102 389174
rect 100186 388938 100422 389174
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 99866 317258 100102 317494
rect 100186 317258 100422 317494
rect 99866 316938 100102 317174
rect 100186 316938 100422 317174
rect 99866 281258 100102 281494
rect 100186 281258 100422 281494
rect 99866 280938 100102 281174
rect 100186 280938 100422 281174
rect 99866 245258 100102 245494
rect 100186 245258 100422 245494
rect 99866 244938 100102 245174
rect 100186 244938 100422 245174
rect 99866 209258 100102 209494
rect 100186 209258 100422 209494
rect 99866 208938 100102 209174
rect 100186 208938 100422 209174
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 124706 486098 124942 486334
rect 125026 486098 125262 486334
rect 124706 485778 124942 486014
rect 125026 485778 125262 486014
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 124706 414098 124942 414334
rect 125026 414098 125262 414334
rect 124706 413778 124942 414014
rect 125026 413778 125262 414014
rect 124706 378098 124942 378334
rect 125026 378098 125262 378334
rect 124706 377778 124942 378014
rect 125026 377778 125262 378014
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 128426 489818 128662 490054
rect 128746 489818 128982 490054
rect 128426 489498 128662 489734
rect 128746 489498 128982 489734
rect 128426 453818 128662 454054
rect 128746 453818 128982 454054
rect 128426 453498 128662 453734
rect 128746 453498 128982 453734
rect 128426 417818 128662 418054
rect 128746 417818 128982 418054
rect 128426 417498 128662 417734
rect 128746 417498 128982 417734
rect 128426 381818 128662 382054
rect 128746 381818 128982 382054
rect 128426 381498 128662 381734
rect 128746 381498 128982 381734
rect 128426 345818 128662 346054
rect 128746 345818 128982 346054
rect 128426 345498 128662 345734
rect 128746 345498 128982 345734
rect 128426 309818 128662 310054
rect 128746 309818 128982 310054
rect 128426 309498 128662 309734
rect 128746 309498 128982 309734
rect 128426 273818 128662 274054
rect 128746 273818 128982 274054
rect 128426 273498 128662 273734
rect 128746 273498 128982 273734
rect 128426 237818 128662 238054
rect 128746 237818 128982 238054
rect 128426 237498 128662 237734
rect 128746 237498 128982 237734
rect 128426 201818 128662 202054
rect 128746 201818 128982 202054
rect 128426 201498 128662 201734
rect 128746 201498 128982 201734
rect 132146 493538 132382 493774
rect 132466 493538 132702 493774
rect 132146 493218 132382 493454
rect 132466 493218 132702 493454
rect 132146 457538 132382 457774
rect 132466 457538 132702 457774
rect 132146 457218 132382 457454
rect 132466 457218 132702 457454
rect 132146 421538 132382 421774
rect 132466 421538 132702 421774
rect 132146 421218 132382 421454
rect 132466 421218 132702 421454
rect 132146 385538 132382 385774
rect 132466 385538 132702 385774
rect 132146 385218 132382 385454
rect 132466 385218 132702 385454
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 135866 497258 136102 497494
rect 136186 497258 136422 497494
rect 135866 496938 136102 497174
rect 136186 496938 136422 497174
rect 135866 461258 136102 461494
rect 136186 461258 136422 461494
rect 135866 460938 136102 461174
rect 136186 460938 136422 461174
rect 135866 425258 136102 425494
rect 136186 425258 136422 425494
rect 135866 424938 136102 425174
rect 136186 424938 136422 425174
rect 135866 389258 136102 389494
rect 136186 389258 136422 389494
rect 135866 388938 136102 389174
rect 136186 388938 136422 389174
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 160706 486098 160942 486334
rect 161026 486098 161262 486334
rect 160706 485778 160942 486014
rect 161026 485778 161262 486014
rect 160706 450098 160942 450334
rect 161026 450098 161262 450334
rect 160706 449778 160942 450014
rect 161026 449778 161262 450014
rect 160706 414098 160942 414334
rect 161026 414098 161262 414334
rect 160706 413778 160942 414014
rect 161026 413778 161262 414014
rect 160706 378098 160942 378334
rect 161026 378098 161262 378334
rect 160706 377778 160942 378014
rect 161026 377778 161262 378014
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 20328 186938 20564 187174
rect 20328 186618 20564 186854
rect 156056 186938 156292 187174
rect 156056 186618 156292 186854
rect 21008 183218 21244 183454
rect 21008 182898 21244 183134
rect 155376 183218 155612 183454
rect 155376 182898 155612 183134
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 20328 150938 20564 151174
rect 20328 150618 20564 150854
rect 156056 150938 156292 151174
rect 156056 150618 156292 150854
rect 21008 147218 21244 147454
rect 21008 146898 21244 147134
rect 155376 147218 155612 147454
rect 155376 146898 155612 147134
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 20328 114938 20564 115174
rect 20328 114618 20564 114854
rect 156056 114938 156292 115174
rect 156056 114618 156292 114854
rect 21008 111101 21244 111337
rect 155376 111101 155612 111337
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 20328 78938 20564 79174
rect 20328 78618 20564 78854
rect 156056 78938 156292 79174
rect 156056 78618 156292 78854
rect 21008 75218 21244 75454
rect 21008 74898 21244 75134
rect 155376 75218 155612 75454
rect 155376 74898 155612 75134
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 20328 42938 20564 43174
rect 20328 42618 20564 42854
rect 156056 42938 156292 43174
rect 156056 42618 156292 42854
rect 21008 39218 21244 39454
rect 21008 38898 21244 39134
rect 155376 39218 155612 39454
rect 155376 38898 155612 39134
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 17787 52942 18023
rect 53026 17787 53262 18023
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 88706 17787 88942 18023
rect 89026 17787 89262 18023
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 124706 17787 124942 18023
rect 125026 17787 125262 18023
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 164426 597818 164662 598054
rect 164746 597818 164982 598054
rect 164426 597498 164662 597734
rect 164746 597498 164982 597734
rect 164426 561818 164662 562054
rect 164746 561818 164982 562054
rect 164426 561498 164662 561734
rect 164746 561498 164982 561734
rect 164426 525818 164662 526054
rect 164746 525818 164982 526054
rect 164426 525498 164662 525734
rect 164746 525498 164982 525734
rect 164426 489818 164662 490054
rect 164746 489818 164982 490054
rect 164426 489498 164662 489734
rect 164746 489498 164982 489734
rect 164426 453818 164662 454054
rect 164746 453818 164982 454054
rect 164426 453498 164662 453734
rect 164746 453498 164982 453734
rect 164426 417818 164662 418054
rect 164746 417818 164982 418054
rect 164426 417498 164662 417734
rect 164746 417498 164982 417734
rect 164426 381818 164662 382054
rect 164746 381818 164982 382054
rect 164426 381498 164662 381734
rect 164746 381498 164982 381734
rect 164426 345818 164662 346054
rect 164746 345818 164982 346054
rect 164426 345498 164662 345734
rect 164746 345498 164982 345734
rect 164426 309818 164662 310054
rect 164746 309818 164982 310054
rect 164426 309498 164662 309734
rect 164746 309498 164982 309734
rect 164426 273818 164662 274054
rect 164746 273818 164982 274054
rect 164426 273498 164662 273734
rect 164746 273498 164982 273734
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 164426 129818 164662 130054
rect 164746 129818 164982 130054
rect 164426 129498 164662 129734
rect 164746 129498 164982 129734
rect 164426 93818 164662 94054
rect 164746 93818 164982 94054
rect 164426 93498 164662 93734
rect 164746 93498 164982 93734
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 168146 601538 168382 601774
rect 168466 601538 168702 601774
rect 168146 601218 168382 601454
rect 168466 601218 168702 601454
rect 168146 565538 168382 565774
rect 168466 565538 168702 565774
rect 168146 565218 168382 565454
rect 168466 565218 168702 565454
rect 168146 529538 168382 529774
rect 168466 529538 168702 529774
rect 168146 529218 168382 529454
rect 168466 529218 168702 529454
rect 168146 493538 168382 493774
rect 168466 493538 168702 493774
rect 168146 493218 168382 493454
rect 168466 493218 168702 493454
rect 168146 457538 168382 457774
rect 168466 457538 168702 457774
rect 168146 457218 168382 457454
rect 168466 457218 168702 457454
rect 168146 421538 168382 421774
rect 168466 421538 168702 421774
rect 168146 421218 168382 421454
rect 168466 421218 168702 421454
rect 168146 385538 168382 385774
rect 168466 385538 168702 385774
rect 168146 385218 168382 385454
rect 168466 385218 168702 385454
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 171866 605258 172102 605494
rect 172186 605258 172422 605494
rect 171866 604938 172102 605174
rect 172186 604938 172422 605174
rect 171866 569258 172102 569494
rect 172186 569258 172422 569494
rect 171866 568938 172102 569174
rect 172186 568938 172422 569174
rect 171866 533258 172102 533494
rect 172186 533258 172422 533494
rect 171866 532938 172102 533174
rect 172186 532938 172422 533174
rect 171866 497258 172102 497494
rect 172186 497258 172422 497494
rect 171866 496938 172102 497174
rect 172186 496938 172422 497174
rect 171866 461258 172102 461494
rect 172186 461258 172422 461494
rect 171866 460938 172102 461174
rect 172186 460938 172422 461174
rect 171866 425258 172102 425494
rect 172186 425258 172422 425494
rect 171866 424938 172102 425174
rect 172186 424938 172422 425174
rect 171866 389258 172102 389494
rect 172186 389258 172422 389494
rect 171866 388938 172102 389174
rect 172186 388938 172422 389174
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 196706 630098 196942 630334
rect 197026 630098 197262 630334
rect 196706 629778 196942 630014
rect 197026 629778 197262 630014
rect 196706 594098 196942 594334
rect 197026 594098 197262 594334
rect 196706 593778 196942 594014
rect 197026 593778 197262 594014
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 196706 486098 196942 486334
rect 197026 486098 197262 486334
rect 196706 485778 196942 486014
rect 197026 485778 197262 486014
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 200426 597818 200662 598054
rect 200746 597818 200982 598054
rect 200426 597498 200662 597734
rect 200746 597498 200982 597734
rect 200426 561818 200662 562054
rect 200746 561818 200982 562054
rect 200426 561498 200662 561734
rect 200746 561498 200982 561734
rect 200426 525818 200662 526054
rect 200746 525818 200982 526054
rect 200426 525498 200662 525734
rect 200746 525498 200982 525734
rect 200426 489818 200662 490054
rect 200746 489818 200982 490054
rect 200426 489498 200662 489734
rect 200746 489498 200982 489734
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 194250 435218 194486 435454
rect 194250 434898 194486 435134
rect 196706 414098 196942 414334
rect 197026 414098 197262 414334
rect 196706 413778 196942 414014
rect 197026 413778 197262 414014
rect 194250 399218 194486 399454
rect 194250 398898 194486 399134
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 194250 363218 194486 363454
rect 194250 362898 194486 363134
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 194250 327218 194486 327454
rect 194250 326898 194486 327134
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 194250 291218 194486 291454
rect 194250 290898 194486 291134
rect 196706 270098 196942 270334
rect 197026 270098 197262 270334
rect 196706 269778 196942 270014
rect 197026 269778 197262 270014
rect 194250 255218 194486 255454
rect 194250 254898 194486 255134
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 196706 198098 196942 198334
rect 197026 198098 197262 198334
rect 196706 197778 196942 198014
rect 197026 197778 197262 198014
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 453818 200662 454054
rect 200746 453818 200982 454054
rect 200426 453498 200662 453734
rect 200746 453498 200982 453734
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 204250 651218 204486 651454
rect 204250 650898 204486 651134
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 204250 615218 204486 615454
rect 204250 614898 204486 615134
rect 207866 605258 208102 605494
rect 208186 605258 208422 605494
rect 207866 604938 208102 605174
rect 208186 604938 208422 605174
rect 204250 579218 204486 579454
rect 204250 578898 204486 579134
rect 207866 569258 208102 569494
rect 208186 569258 208422 569494
rect 207866 568938 208102 569174
rect 208186 568938 208422 569174
rect 204250 543218 204486 543454
rect 204250 542898 204486 543134
rect 207866 533258 208102 533494
rect 208186 533258 208422 533494
rect 207866 532938 208102 533174
rect 208186 532938 208422 533174
rect 204250 507218 204486 507454
rect 204250 506898 204486 507134
rect 204146 493538 204382 493774
rect 204466 493538 204702 493774
rect 204146 493218 204382 493454
rect 204466 493218 204702 493454
rect 204146 457538 204382 457774
rect 204466 457538 204702 457774
rect 204146 457218 204382 457454
rect 204466 457218 204702 457454
rect 200426 417818 200662 418054
rect 200746 417818 200982 418054
rect 200426 417498 200662 417734
rect 200746 417498 200982 417734
rect 200426 381818 200662 382054
rect 200746 381818 200982 382054
rect 200426 381498 200662 381734
rect 200746 381498 200982 381734
rect 200426 345818 200662 346054
rect 200746 345818 200982 346054
rect 200426 345498 200662 345734
rect 200746 345498 200982 345734
rect 200426 309818 200662 310054
rect 200746 309818 200982 310054
rect 200426 309498 200662 309734
rect 200746 309498 200982 309734
rect 200426 273818 200662 274054
rect 200746 273818 200982 274054
rect 200426 273498 200662 273734
rect 200746 273498 200982 273734
rect 200426 237818 200662 238054
rect 200746 237818 200982 238054
rect 200426 237498 200662 237734
rect 200746 237498 200982 237734
rect 200426 201818 200662 202054
rect 200746 201818 200982 202054
rect 200426 201498 200662 201734
rect 200746 201498 200982 201734
rect 200426 165818 200662 166054
rect 200746 165818 200982 166054
rect 200426 165498 200662 165734
rect 200746 165498 200982 165734
rect 200426 129818 200662 130054
rect 200746 129818 200982 130054
rect 200426 129498 200662 129734
rect 200746 129498 200982 129734
rect 200426 93818 200662 94054
rect 200746 93818 200982 94054
rect 200426 93498 200662 93734
rect 200746 93498 200982 93734
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 421538 204382 421774
rect 204466 421538 204702 421774
rect 204146 421218 204382 421454
rect 204466 421218 204702 421454
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 204146 277538 204382 277774
rect 204466 277538 204702 277774
rect 204146 277218 204382 277454
rect 204466 277218 204702 277454
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 204146 205538 204382 205774
rect 204466 205538 204702 205774
rect 204146 205218 204382 205454
rect 204466 205218 204702 205454
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 497258 208102 497494
rect 208186 497258 208422 497494
rect 207866 496938 208102 497174
rect 208186 496938 208422 497174
rect 207866 461258 208102 461494
rect 208186 461258 208422 461494
rect 207866 460938 208102 461174
rect 208186 460938 208422 461174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 219610 654938 219846 655174
rect 219610 654618 219846 654854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 219610 618938 219846 619174
rect 219610 618618 219846 618854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 219610 582938 219846 583174
rect 219610 582618 219846 582854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 219610 546938 219846 547174
rect 219610 546618 219846 546854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 219610 510938 219846 511174
rect 219610 510618 219846 510854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 209610 438938 209846 439174
rect 209610 438618 209846 438854
rect 207866 425258 208102 425494
rect 208186 425258 208422 425494
rect 207866 424938 208102 425174
rect 208186 424938 208422 425174
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 209610 402938 209846 403174
rect 209610 402618 209846 402854
rect 207866 389258 208102 389494
rect 208186 389258 208422 389494
rect 207866 388938 208102 389174
rect 208186 388938 208422 389174
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 209610 366938 209846 367174
rect 209610 366618 209846 366854
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 209610 330938 209846 331174
rect 209610 330618 209846 330854
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 209610 294938 209846 295174
rect 209610 294618 209846 294854
rect 207866 281258 208102 281494
rect 208186 281258 208422 281494
rect 207866 280938 208102 281174
rect 208186 280938 208422 281174
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 209610 258938 209846 259174
rect 209610 258618 209846 258854
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 207866 209258 208102 209494
rect 208186 209258 208422 209494
rect 207866 208938 208102 209174
rect 208186 208938 208422 209174
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 224970 435218 225206 435454
rect 224970 434898 225206 435134
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 224970 399218 225206 399454
rect 224970 398898 225206 399134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 224970 363218 225206 363454
rect 224970 362898 225206 363134
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 224970 327218 225206 327454
rect 224970 326898 225206 327134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 224970 291218 225206 291454
rect 224970 290898 225206 291134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 224970 255218 225206 255454
rect 224970 254898 225206 255134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 234970 651218 235206 651454
rect 234970 650898 235206 651134
rect 232706 630098 232942 630334
rect 233026 630098 233262 630334
rect 232706 629778 232942 630014
rect 233026 629778 233262 630014
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 234970 615218 235206 615454
rect 234970 614898 235206 615134
rect 232706 594098 232942 594334
rect 233026 594098 233262 594334
rect 232706 593778 232942 594014
rect 233026 593778 233262 594014
rect 236426 597818 236662 598054
rect 236746 597818 236982 598054
rect 236426 597498 236662 597734
rect 236746 597498 236982 597734
rect 234970 579218 235206 579454
rect 234970 578898 235206 579134
rect 232706 558098 232942 558334
rect 233026 558098 233262 558334
rect 232706 557778 232942 558014
rect 233026 557778 233262 558014
rect 236426 561818 236662 562054
rect 236746 561818 236982 562054
rect 236426 561498 236662 561734
rect 236746 561498 236982 561734
rect 234970 543218 235206 543454
rect 234970 542898 235206 543134
rect 232706 522098 232942 522334
rect 233026 522098 233262 522334
rect 232706 521778 232942 522014
rect 233026 521778 233262 522014
rect 236426 525818 236662 526054
rect 236746 525818 236982 526054
rect 236426 525498 236662 525734
rect 236746 525498 236982 525734
rect 234970 507218 235206 507454
rect 234970 506898 235206 507134
rect 232706 486098 232942 486334
rect 233026 486098 233262 486334
rect 232706 485778 232942 486014
rect 233026 485778 233262 486014
rect 232706 450098 232942 450334
rect 233026 450098 233262 450334
rect 232706 449778 232942 450014
rect 233026 449778 233262 450014
rect 232706 414098 232942 414334
rect 233026 414098 233262 414334
rect 232706 413778 232942 414014
rect 233026 413778 233262 414014
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 236426 489818 236662 490054
rect 236746 489818 236982 490054
rect 236426 489498 236662 489734
rect 236746 489498 236982 489734
rect 236426 453818 236662 454054
rect 236746 453818 236982 454054
rect 236426 453498 236662 453734
rect 236746 453498 236982 453734
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 250330 654938 250566 655174
rect 250330 654618 250566 654854
rect 281050 654938 281286 655174
rect 281050 654618 281286 654854
rect 311770 654938 312006 655174
rect 311770 654618 312006 654854
rect 265690 651218 265926 651454
rect 265690 650898 265926 651134
rect 296410 651218 296646 651454
rect 296410 650898 296646 651134
rect 327130 651218 327366 651454
rect 327130 650898 327366 651134
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 250330 618938 250566 619174
rect 250330 618618 250566 618854
rect 281050 618938 281286 619174
rect 281050 618618 281286 618854
rect 311770 618938 312006 619174
rect 311770 618618 312006 618854
rect 265690 615218 265926 615454
rect 265690 614898 265926 615134
rect 296410 615218 296646 615454
rect 296410 614898 296646 615134
rect 327130 615218 327366 615454
rect 327130 614898 327366 615134
rect 240146 601538 240382 601774
rect 240466 601538 240702 601774
rect 240146 601218 240382 601454
rect 240466 601218 240702 601454
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 250330 582938 250566 583174
rect 250330 582618 250566 582854
rect 281050 582938 281286 583174
rect 281050 582618 281286 582854
rect 311770 582938 312006 583174
rect 311770 582618 312006 582854
rect 265690 579218 265926 579454
rect 265690 578898 265926 579134
rect 296410 579218 296646 579454
rect 296410 578898 296646 579134
rect 327130 579218 327366 579454
rect 327130 578898 327366 579134
rect 240146 565538 240382 565774
rect 240466 565538 240702 565774
rect 240146 565218 240382 565454
rect 240466 565218 240702 565454
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 250330 546938 250566 547174
rect 250330 546618 250566 546854
rect 281050 546938 281286 547174
rect 281050 546618 281286 546854
rect 311770 546938 312006 547174
rect 311770 546618 312006 546854
rect 265690 543218 265926 543454
rect 265690 542898 265926 543134
rect 296410 543218 296646 543454
rect 296410 542898 296646 543134
rect 327130 543218 327366 543454
rect 327130 542898 327366 543134
rect 240146 529538 240382 529774
rect 240466 529538 240702 529774
rect 240146 529218 240382 529454
rect 240466 529218 240702 529454
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 250330 510938 250566 511174
rect 250330 510618 250566 510854
rect 281050 510938 281286 511174
rect 281050 510618 281286 510854
rect 311770 510938 312006 511174
rect 311770 510618 312006 510854
rect 265690 507218 265926 507454
rect 265690 506898 265926 507134
rect 296410 507218 296646 507454
rect 296410 506898 296646 507134
rect 327130 507218 327366 507454
rect 327130 506898 327366 507134
rect 240146 493538 240382 493774
rect 240466 493538 240702 493774
rect 240146 493218 240382 493454
rect 240466 493218 240702 493454
rect 240146 457538 240382 457774
rect 240466 457538 240702 457774
rect 240146 457218 240382 457454
rect 240466 457218 240702 457454
rect 243866 497258 244102 497494
rect 244186 497258 244422 497494
rect 243866 496938 244102 497174
rect 244186 496938 244422 497174
rect 243866 461258 244102 461494
rect 244186 461258 244422 461494
rect 243866 460938 244102 461174
rect 244186 460938 244422 461174
rect 240330 438938 240566 439174
rect 240330 438618 240566 438854
rect 236426 417818 236662 418054
rect 236746 417818 236982 418054
rect 236426 417498 236662 417734
rect 236746 417498 236982 417734
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 243866 425258 244102 425494
rect 244186 425258 244422 425494
rect 243866 424938 244102 425174
rect 244186 424938 244422 425174
rect 240330 402938 240566 403174
rect 240330 402618 240566 402854
rect 236426 381818 236662 382054
rect 236746 381818 236982 382054
rect 236426 381498 236662 381734
rect 236746 381498 236982 381734
rect 243866 389258 244102 389494
rect 244186 389258 244422 389494
rect 243866 388938 244102 389174
rect 244186 388938 244422 389174
rect 240330 366938 240566 367174
rect 240330 366618 240566 366854
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 243866 353258 244102 353494
rect 244186 353258 244422 353494
rect 243866 352938 244102 353174
rect 244186 352938 244422 353174
rect 240330 330938 240566 331174
rect 240330 330618 240566 330854
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 243866 317258 244102 317494
rect 244186 317258 244422 317494
rect 243866 316938 244102 317174
rect 244186 316938 244422 317174
rect 240330 294938 240566 295174
rect 240330 294618 240566 294854
rect 236426 273818 236662 274054
rect 236746 273818 236982 274054
rect 236426 273498 236662 273734
rect 236746 273498 236982 273734
rect 243866 281258 244102 281494
rect 244186 281258 244422 281494
rect 243866 280938 244102 281174
rect 244186 280938 244422 281174
rect 240330 258938 240566 259174
rect 240330 258618 240566 258854
rect 236426 237818 236662 238054
rect 236746 237818 236982 238054
rect 236426 237498 236662 237734
rect 236746 237498 236982 237734
rect 236426 201818 236662 202054
rect 236746 201818 236982 202054
rect 236426 201498 236662 201734
rect 236746 201498 236982 201734
rect 236426 165818 236662 166054
rect 236746 165818 236982 166054
rect 236426 165498 236662 165734
rect 236746 165498 236982 165734
rect 236426 129818 236662 130054
rect 236746 129818 236982 130054
rect 236426 129498 236662 129734
rect 236746 129498 236982 129734
rect 240146 241538 240382 241774
rect 240466 241538 240702 241774
rect 240146 241218 240382 241454
rect 240466 241218 240702 241454
rect 240146 205538 240382 205774
rect 240466 205538 240702 205774
rect 240146 205218 240382 205454
rect 240466 205218 240702 205454
rect 240146 169538 240382 169774
rect 240466 169538 240702 169774
rect 240146 169218 240382 169454
rect 240466 169218 240702 169454
rect 240146 133538 240382 133774
rect 240466 133538 240702 133774
rect 240146 133218 240382 133454
rect 240466 133218 240702 133454
rect 243866 245258 244102 245494
rect 244186 245258 244422 245494
rect 243866 244938 244102 245174
rect 244186 244938 244422 245174
rect 243866 209258 244102 209494
rect 244186 209258 244422 209494
rect 243866 208938 244102 209174
rect 244186 208938 244422 209174
rect 243866 173258 244102 173494
rect 244186 173258 244422 173494
rect 243866 172938 244102 173174
rect 244186 172938 244422 173174
rect 243866 137258 244102 137494
rect 244186 137258 244422 137494
rect 243866 136938 244102 137174
rect 244186 136938 244422 137174
rect 272426 489818 272662 490054
rect 272746 489818 272982 490054
rect 272426 489498 272662 489734
rect 272746 489498 272982 489734
rect 272426 453818 272662 454054
rect 272746 453818 272982 454054
rect 272426 453498 272662 453734
rect 272746 453498 272982 453734
rect 276146 493538 276382 493774
rect 276466 493538 276702 493774
rect 276146 493218 276382 493454
rect 276466 493218 276702 493454
rect 276146 457538 276382 457774
rect 276466 457538 276702 457774
rect 276146 457218 276382 457454
rect 276466 457218 276702 457454
rect 279866 497258 280102 497494
rect 280186 497258 280422 497494
rect 279866 496938 280102 497174
rect 280186 496938 280422 497174
rect 279866 461258 280102 461494
rect 280186 461258 280422 461494
rect 279866 460938 280102 461174
rect 280186 460938 280422 461174
rect 308426 489818 308662 490054
rect 308746 489818 308982 490054
rect 308426 489498 308662 489734
rect 308746 489498 308982 489734
rect 308426 453818 308662 454054
rect 308746 453818 308982 454054
rect 308426 453498 308662 453734
rect 308746 453498 308982 453734
rect 312146 493538 312382 493774
rect 312466 493538 312702 493774
rect 312146 493218 312382 493454
rect 312466 493218 312702 493454
rect 312146 457538 312382 457774
rect 312466 457538 312702 457774
rect 312146 457218 312382 457454
rect 312466 457218 312702 457454
rect 315866 497258 316102 497494
rect 316186 497258 316422 497494
rect 315866 496938 316102 497174
rect 316186 496938 316422 497174
rect 315866 461258 316102 461494
rect 316186 461258 316422 461494
rect 315866 460938 316102 461174
rect 316186 460938 316422 461174
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 342490 654938 342726 655174
rect 342490 654618 342726 654854
rect 340706 630098 340942 630334
rect 341026 630098 341262 630334
rect 340706 629778 340942 630014
rect 341026 629778 341262 630014
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 342490 618938 342726 619174
rect 342490 618618 342726 618854
rect 340706 594098 340942 594334
rect 341026 594098 341262 594334
rect 340706 593778 340942 594014
rect 341026 593778 341262 594014
rect 344426 597818 344662 598054
rect 344746 597818 344982 598054
rect 344426 597498 344662 597734
rect 344746 597498 344982 597734
rect 342490 582938 342726 583174
rect 342490 582618 342726 582854
rect 340706 558098 340942 558334
rect 341026 558098 341262 558334
rect 340706 557778 340942 558014
rect 341026 557778 341262 558014
rect 344426 561818 344662 562054
rect 344746 561818 344982 562054
rect 344426 561498 344662 561734
rect 344746 561498 344982 561734
rect 342490 546938 342726 547174
rect 342490 546618 342726 546854
rect 340706 522098 340942 522334
rect 341026 522098 341262 522334
rect 340706 521778 340942 522014
rect 341026 521778 341262 522014
rect 344426 525818 344662 526054
rect 344746 525818 344982 526054
rect 344426 525498 344662 525734
rect 344746 525498 344982 525734
rect 342490 510938 342726 511174
rect 342490 510618 342726 510854
rect 340706 486098 340942 486334
rect 341026 486098 341262 486334
rect 340706 485778 340942 486014
rect 341026 485778 341262 486014
rect 344426 489818 344662 490054
rect 344746 489818 344982 490054
rect 344426 489498 344662 489734
rect 344746 489498 344982 489734
rect 344426 453818 344662 454054
rect 344746 453818 344982 454054
rect 344426 453498 344662 453734
rect 344746 453498 344982 453734
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 348146 601538 348382 601774
rect 348466 601538 348702 601774
rect 348146 601218 348382 601454
rect 348466 601218 348702 601454
rect 348146 565538 348382 565774
rect 348466 565538 348702 565774
rect 348146 565218 348382 565454
rect 348466 565218 348702 565454
rect 348146 529538 348382 529774
rect 348466 529538 348702 529774
rect 348146 529218 348382 529454
rect 348466 529218 348702 529454
rect 348146 493538 348382 493774
rect 348466 493538 348702 493774
rect 348146 493218 348382 493454
rect 348466 493218 348702 493454
rect 348146 457538 348382 457774
rect 348466 457538 348702 457774
rect 348146 457218 348382 457454
rect 348466 457218 348702 457454
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 357850 651218 358086 651454
rect 357850 650898 358086 651134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 357850 615218 358086 615454
rect 357850 614898 358086 615134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 351866 605258 352102 605494
rect 352186 605258 352422 605494
rect 351866 604938 352102 605174
rect 352186 604938 352422 605174
rect 357850 579218 358086 579454
rect 357850 578898 358086 579134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 351866 569258 352102 569494
rect 352186 569258 352422 569494
rect 351866 568938 352102 569174
rect 352186 568938 352422 569174
rect 357850 543218 358086 543454
rect 357850 542898 358086 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 351866 533258 352102 533494
rect 352186 533258 352422 533494
rect 351866 532938 352102 533174
rect 352186 532938 352422 533174
rect 357850 507218 358086 507454
rect 357850 506898 358086 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 351866 497258 352102 497494
rect 352186 497258 352422 497494
rect 351866 496938 352102 497174
rect 352186 496938 352422 497174
rect 351866 461258 352102 461494
rect 352186 461258 352422 461494
rect 351866 460938 352102 461174
rect 352186 460938 352422 461174
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 373210 654938 373446 655174
rect 373210 654618 373446 654854
rect 373210 618938 373446 619174
rect 373210 618618 373446 618854
rect 373210 582938 373446 583174
rect 373210 582618 373446 582854
rect 373210 546938 373446 547174
rect 373210 546618 373446 546854
rect 373210 510938 373446 511174
rect 373210 510618 373446 510854
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 271050 438938 271286 439174
rect 271050 438618 271286 438854
rect 301770 438938 302006 439174
rect 301770 438618 302006 438854
rect 332490 438938 332726 439174
rect 332490 438618 332726 438854
rect 363210 438938 363446 439174
rect 363210 438618 363446 438854
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 255690 435218 255926 435454
rect 255690 434898 255926 435134
rect 286410 435218 286646 435454
rect 286410 434898 286646 435134
rect 317130 435218 317366 435454
rect 317130 434898 317366 435134
rect 347850 435218 348086 435454
rect 347850 434898 348086 435134
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 271050 402938 271286 403174
rect 271050 402618 271286 402854
rect 301770 402938 302006 403174
rect 301770 402618 302006 402854
rect 332490 402938 332726 403174
rect 332490 402618 332726 402854
rect 363210 402938 363446 403174
rect 363210 402618 363446 402854
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 255690 399218 255926 399454
rect 255690 398898 255926 399134
rect 286410 399218 286646 399454
rect 286410 398898 286646 399134
rect 317130 399218 317366 399454
rect 317130 398898 317366 399134
rect 347850 399218 348086 399454
rect 347850 398898 348086 399134
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 271050 366938 271286 367174
rect 271050 366618 271286 366854
rect 301770 366938 302006 367174
rect 301770 366618 302006 366854
rect 332490 366938 332726 367174
rect 332490 366618 332726 366854
rect 363210 366938 363446 367174
rect 363210 366618 363446 366854
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 255690 363218 255926 363454
rect 255690 362898 255926 363134
rect 286410 363218 286646 363454
rect 286410 362898 286646 363134
rect 317130 363218 317366 363454
rect 317130 362898 317366 363134
rect 347850 363218 348086 363454
rect 347850 362898 348086 363134
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 271050 330938 271286 331174
rect 271050 330618 271286 330854
rect 301770 330938 302006 331174
rect 301770 330618 302006 330854
rect 332490 330938 332726 331174
rect 332490 330618 332726 330854
rect 363210 330938 363446 331174
rect 363210 330618 363446 330854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 255690 327218 255926 327454
rect 255690 326898 255926 327134
rect 286410 327218 286646 327454
rect 286410 326898 286646 327134
rect 317130 327218 317366 327454
rect 317130 326898 317366 327134
rect 347850 327218 348086 327454
rect 347850 326898 348086 327134
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 271050 294938 271286 295174
rect 271050 294618 271286 294854
rect 301770 294938 302006 295174
rect 301770 294618 302006 294854
rect 332490 294938 332726 295174
rect 332490 294618 332726 294854
rect 363210 294938 363446 295174
rect 363210 294618 363446 294854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 255690 291218 255926 291454
rect 255690 290898 255926 291134
rect 286410 291218 286646 291454
rect 286410 290898 286646 291134
rect 317130 291218 317366 291454
rect 317130 290898 317366 291134
rect 347850 291218 348086 291454
rect 347850 290898 348086 291134
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 271050 258938 271286 259174
rect 271050 258618 271286 258854
rect 301770 258938 302006 259174
rect 301770 258618 302006 258854
rect 332490 258938 332726 259174
rect 332490 258618 332726 258854
rect 363210 258938 363446 259174
rect 363210 258618 363446 258854
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 255690 255218 255926 255454
rect 255690 254898 255926 255134
rect 286410 255218 286646 255454
rect 286410 254898 286646 255134
rect 317130 255218 317366 255454
rect 317130 254898 317366 255134
rect 347850 255218 348086 255454
rect 347850 254898 348086 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 268706 234098 268942 234334
rect 269026 234098 269262 234334
rect 268706 233778 268942 234014
rect 269026 233778 269262 234014
rect 268706 198098 268942 198334
rect 269026 198098 269262 198334
rect 268706 197778 268942 198014
rect 269026 197778 269262 198014
rect 268706 162098 268942 162334
rect 269026 162098 269262 162334
rect 268706 161778 268942 162014
rect 269026 161778 269262 162014
rect 268706 126098 268942 126334
rect 269026 126098 269262 126334
rect 268706 125778 268942 126014
rect 269026 125778 269262 126014
rect 272426 237818 272662 238054
rect 272746 237818 272982 238054
rect 272426 237498 272662 237734
rect 272746 237498 272982 237734
rect 272426 201818 272662 202054
rect 272746 201818 272982 202054
rect 272426 201498 272662 201734
rect 272746 201498 272982 201734
rect 272426 165818 272662 166054
rect 272746 165818 272982 166054
rect 272426 165498 272662 165734
rect 272746 165498 272982 165734
rect 272426 129818 272662 130054
rect 272746 129818 272982 130054
rect 272426 129498 272662 129734
rect 272746 129498 272982 129734
rect 276146 241538 276382 241774
rect 276466 241538 276702 241774
rect 276146 241218 276382 241454
rect 276466 241218 276702 241454
rect 276146 205538 276382 205774
rect 276466 205538 276702 205774
rect 276146 205218 276382 205454
rect 276466 205218 276702 205454
rect 276146 169538 276382 169774
rect 276466 169538 276702 169774
rect 276146 169218 276382 169454
rect 276466 169218 276702 169454
rect 276146 133538 276382 133774
rect 276466 133538 276702 133774
rect 276146 133218 276382 133454
rect 276466 133218 276702 133454
rect 279866 245258 280102 245494
rect 280186 245258 280422 245494
rect 279866 244938 280102 245174
rect 280186 244938 280422 245174
rect 279866 209258 280102 209494
rect 280186 209258 280422 209494
rect 279866 208938 280102 209174
rect 280186 208938 280422 209174
rect 279866 173258 280102 173494
rect 280186 173258 280422 173494
rect 279866 172938 280102 173174
rect 280186 172938 280422 173174
rect 279866 137258 280102 137494
rect 280186 137258 280422 137494
rect 279866 136938 280102 137174
rect 280186 136938 280422 137174
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 308426 237818 308662 238054
rect 308746 237818 308982 238054
rect 308426 237498 308662 237734
rect 308746 237498 308982 237734
rect 308426 201818 308662 202054
rect 308746 201818 308982 202054
rect 308426 201498 308662 201734
rect 308746 201498 308982 201734
rect 308426 165818 308662 166054
rect 308746 165818 308982 166054
rect 308426 165498 308662 165734
rect 308746 165498 308982 165734
rect 308426 129818 308662 130054
rect 308746 129818 308982 130054
rect 308426 129498 308662 129734
rect 308746 129498 308982 129734
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 340706 234098 340942 234334
rect 341026 234098 341262 234334
rect 340706 233778 340942 234014
rect 341026 233778 341262 234014
rect 340706 198098 340942 198334
rect 341026 198098 341262 198334
rect 340706 197778 340942 198014
rect 341026 197778 341262 198014
rect 340706 162098 340942 162334
rect 341026 162098 341262 162334
rect 340706 161778 340942 162014
rect 341026 161778 341262 162014
rect 340706 126098 340942 126334
rect 341026 126098 341262 126334
rect 340706 125778 340942 126014
rect 341026 125778 341262 126014
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 207866 101258 208102 101494
rect 208186 101258 208422 101494
rect 207866 100938 208102 101174
rect 208186 100938 208422 101174
rect 220328 78938 220564 79174
rect 220328 78618 220564 78854
rect 356056 78938 356292 79174
rect 356056 78618 356292 78854
rect 221008 75218 221244 75454
rect 221008 74898 221244 75134
rect 355376 75218 355612 75454
rect 355376 74898 355612 75134
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 220328 42938 220564 43174
rect 220328 42618 220564 42854
rect 356056 42938 356292 43174
rect 356056 42618 356292 42854
rect 221008 39218 221244 39454
rect 221008 38898 221244 39134
rect 355376 39218 355612 39454
rect 355376 38898 355612 39134
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 17787 232942 18023
rect 233026 17787 233262 18023
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 17787 304942 18023
rect 305026 17787 305262 18023
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 17787 340942 18023
rect 341026 17787 341262 18023
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 378570 435218 378806 435454
rect 378570 434898 378806 435134
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 378570 399218 378806 399454
rect 378570 398898 378806 399134
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 378570 363218 378806 363454
rect 378570 362898 378806 363134
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 378570 327218 378806 327454
rect 378570 326898 378806 327134
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 378570 291218 378806 291454
rect 378570 290898 378806 291134
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 378570 255218 378806 255454
rect 378570 254898 378806 255134
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 420328 654938 420564 655174
rect 420328 654618 420564 654854
rect 556056 654938 556292 655174
rect 556056 654618 556292 654854
rect 421008 651218 421244 651454
rect 421008 650898 421244 651134
rect 555376 651218 555612 651454
rect 555376 650898 555612 651134
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 420328 618938 420564 619174
rect 420328 618618 420564 618854
rect 556056 618938 556292 619174
rect 556056 618618 556292 618854
rect 421008 615218 421244 615454
rect 421008 614898 421244 615134
rect 555376 615218 555612 615454
rect 555376 614898 555612 615134
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 420328 582693 420564 582929
rect 556056 582693 556292 582929
rect 421008 579218 421244 579454
rect 421008 578898 421244 579134
rect 555376 579218 555612 579454
rect 555376 578898 555612 579134
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 420328 546938 420564 547174
rect 420328 546618 420564 546854
rect 556056 546938 556292 547174
rect 556056 546618 556292 546854
rect 421008 543218 421244 543454
rect 421008 542898 421244 543134
rect 555376 543218 555612 543454
rect 555376 542898 555612 543134
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 420328 510938 420564 511174
rect 420328 510618 420564 510854
rect 556056 510938 556292 511174
rect 556056 510618 556292 510854
rect 421008 507218 421244 507454
rect 421008 506898 421244 507134
rect 555376 507218 555612 507454
rect 555376 506898 555612 507134
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 416426 129818 416662 130054
rect 416746 129818 416982 130054
rect 416426 129498 416662 129734
rect 416746 129498 416982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 423866 425258 424102 425494
rect 424186 425258 424422 425494
rect 423866 424938 424102 425174
rect 424186 424938 424422 425174
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 484706 378098 484942 378334
rect 485026 378098 485262 378334
rect 484706 377778 484942 378014
rect 485026 377778 485262 378014
rect 484706 342098 484942 342334
rect 485026 342098 485262 342334
rect 484706 341778 484942 342014
rect 485026 341778 485262 342014
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 484706 234098 484942 234334
rect 485026 234098 485262 234334
rect 484706 233778 484942 234014
rect 485026 233778 485262 234014
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453818 488662 454054
rect 488746 453818 488982 454054
rect 488426 453498 488662 453734
rect 488746 453498 488982 453734
rect 488426 417818 488662 418054
rect 488746 417818 488982 418054
rect 488426 417498 488662 417734
rect 488746 417498 488982 417734
rect 488426 381818 488662 382054
rect 488746 381818 488982 382054
rect 488426 381498 488662 381734
rect 488746 381498 488982 381734
rect 488426 345818 488662 346054
rect 488746 345818 488982 346054
rect 488426 345498 488662 345734
rect 488746 345498 488982 345734
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 488426 237818 488662 238054
rect 488746 237818 488982 238054
rect 488426 237498 488662 237734
rect 488746 237498 488982 237734
rect 488426 201818 488662 202054
rect 488746 201818 488982 202054
rect 488426 201498 488662 201734
rect 488746 201498 488982 201734
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 492146 385538 492382 385774
rect 492466 385538 492702 385774
rect 492146 385218 492382 385454
rect 492466 385218 492702 385454
rect 492146 349538 492382 349774
rect 492466 349538 492702 349774
rect 492146 349218 492382 349454
rect 492466 349218 492702 349454
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 492146 241538 492382 241774
rect 492466 241538 492702 241774
rect 492146 241218 492382 241454
rect 492466 241218 492702 241454
rect 492146 205538 492382 205774
rect 492466 205538 492702 205774
rect 492146 205218 492382 205454
rect 492466 205218 492702 205454
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 495866 245258 496102 245494
rect 496186 245258 496422 245494
rect 495866 244938 496102 245174
rect 496186 244938 496422 245174
rect 495866 209258 496102 209494
rect 496186 209258 496422 209494
rect 495866 208938 496102 209174
rect 496186 208938 496422 209174
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 520706 234098 520942 234334
rect 521026 234098 521262 234334
rect 520706 233778 520942 234014
rect 521026 233778 521262 234014
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 524426 237818 524662 238054
rect 524746 237818 524982 238054
rect 524426 237498 524662 237734
rect 524746 237498 524982 237734
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 528146 241538 528382 241774
rect 528466 241538 528702 241774
rect 528146 241218 528382 241454
rect 528466 241218 528702 241454
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 420328 186938 420564 187174
rect 420328 186618 420564 186854
rect 556056 186938 556292 187174
rect 556056 186618 556292 186854
rect 421008 183218 421244 183454
rect 421008 182898 421244 183134
rect 555376 183218 555612 183454
rect 555376 182898 555612 183134
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 420328 150938 420564 151174
rect 420328 150618 420564 150854
rect 556056 150938 556292 151174
rect 556056 150618 556292 150854
rect 421008 147218 421244 147454
rect 421008 146898 421244 147134
rect 555376 147218 555612 147454
rect 555376 146898 555612 147134
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 420328 114938 420564 115174
rect 420328 114618 420564 114854
rect 556056 114938 556292 115174
rect 556056 114618 556292 114854
rect 421008 111101 421244 111337
rect 555376 111101 555612 111337
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 420328 78938 420564 79174
rect 420328 78618 420564 78854
rect 556056 78938 556292 79174
rect 556056 78618 556292 78854
rect 421008 75218 421244 75454
rect 421008 74898 421244 75134
rect 555376 75218 555612 75454
rect 555376 74898 555612 75134
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 420328 42938 420564 43174
rect 420328 42618 420564 42854
rect 556056 42938 556292 43174
rect 556056 42618 556292 42854
rect 421008 39218 421244 39454
rect 421008 38898 421244 39134
rect 555376 39218 555612 39454
rect 555376 38898 555612 39134
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 484706 17787 484942 18023
rect 485026 17787 485262 18023
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 17787 556942 18023
rect 557026 17787 557262 18023
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 20328 655174
rect 20564 654938 156056 655174
rect 156292 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 219610 655174
rect 219846 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 250330 655174
rect 250566 654938 281050 655174
rect 281286 654938 311770 655174
rect 312006 654938 342490 655174
rect 342726 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 373210 655174
rect 373446 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 420328 655174
rect 420564 654938 556056 655174
rect 556292 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 20328 654854
rect 20564 654618 156056 654854
rect 156292 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 219610 654854
rect 219846 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 250330 654854
rect 250566 654618 281050 654854
rect 281286 654618 311770 654854
rect 312006 654618 342490 654854
rect 342726 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 373210 654854
rect 373446 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 420328 654854
rect 420564 654618 556056 654854
rect 556292 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 21008 651454
rect 21244 651218 155376 651454
rect 155612 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 204250 651454
rect 204486 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 234970 651454
rect 235206 651218 265690 651454
rect 265926 651218 296410 651454
rect 296646 651218 327130 651454
rect 327366 651218 357850 651454
rect 358086 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 421008 651454
rect 421244 651218 555376 651454
rect 555612 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 21008 651134
rect 21244 650898 155376 651134
rect 155612 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 204250 651134
rect 204486 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 234970 651134
rect 235206 650898 265690 651134
rect 265926 650898 296410 651134
rect 296646 650898 327130 651134
rect 327366 650898 357850 651134
rect 358086 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 421008 651134
rect 421244 650898 555376 651134
rect 555612 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 20328 619174
rect 20564 618938 156056 619174
rect 156292 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 219610 619174
rect 219846 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 250330 619174
rect 250566 618938 281050 619174
rect 281286 618938 311770 619174
rect 312006 618938 342490 619174
rect 342726 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 373210 619174
rect 373446 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 420328 619174
rect 420564 618938 556056 619174
rect 556292 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 20328 618854
rect 20564 618618 156056 618854
rect 156292 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 219610 618854
rect 219846 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 250330 618854
rect 250566 618618 281050 618854
rect 281286 618618 311770 618854
rect 312006 618618 342490 618854
rect 342726 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 373210 618854
rect 373446 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 420328 618854
rect 420564 618618 556056 618854
rect 556292 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 21008 615454
rect 21244 615218 155376 615454
rect 155612 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 204250 615454
rect 204486 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 234970 615454
rect 235206 615218 265690 615454
rect 265926 615218 296410 615454
rect 296646 615218 327130 615454
rect 327366 615218 357850 615454
rect 358086 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 421008 615454
rect 421244 615218 555376 615454
rect 555612 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 21008 615134
rect 21244 614898 155376 615134
rect 155612 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 204250 615134
rect 204486 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 234970 615134
rect 235206 614898 265690 615134
rect 265926 614898 296410 615134
rect 296646 614898 327130 615134
rect 327366 614898 357850 615134
rect 358086 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 421008 615134
rect 421244 614898 555376 615134
rect 555612 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 219610 583174
rect 219846 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 250330 583174
rect 250566 582938 281050 583174
rect 281286 582938 311770 583174
rect 312006 582938 342490 583174
rect 342726 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 373210 583174
rect 373446 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582929 592650 582938
rect -8726 582854 20328 582929
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582693 20328 582854
rect 20564 582693 156056 582929
rect 156292 582854 420328 582929
rect 156292 582693 185546 582854
rect 6102 582618 185546 582693
rect 185782 582618 185866 582854
rect 186102 582618 219610 582854
rect 219846 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 250330 582854
rect 250566 582618 281050 582854
rect 281286 582618 311770 582854
rect 312006 582618 342490 582854
rect 342726 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 373210 582854
rect 373446 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582693 420328 582854
rect 420564 582693 556056 582929
rect 556292 582854 592650 582929
rect 556292 582693 581546 582854
rect 402102 582618 581546 582693
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 21008 579454
rect 21244 579218 155376 579454
rect 155612 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 204250 579454
rect 204486 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 234970 579454
rect 235206 579218 265690 579454
rect 265926 579218 296410 579454
rect 296646 579218 327130 579454
rect 327366 579218 357850 579454
rect 358086 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 421008 579454
rect 421244 579218 555376 579454
rect 555612 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 21008 579134
rect 21244 578898 155376 579134
rect 155612 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 204250 579134
rect 204486 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 234970 579134
rect 235206 578898 265690 579134
rect 265926 578898 296410 579134
rect 296646 578898 327130 579134
rect 327366 578898 357850 579134
rect 358086 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 421008 579134
rect 421244 578898 555376 579134
rect 555612 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 20328 547174
rect 20564 546938 156056 547174
rect 156292 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 219610 547174
rect 219846 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 250330 547174
rect 250566 546938 281050 547174
rect 281286 546938 311770 547174
rect 312006 546938 342490 547174
rect 342726 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 373210 547174
rect 373446 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 420328 547174
rect 420564 546938 556056 547174
rect 556292 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 20328 546854
rect 20564 546618 156056 546854
rect 156292 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 219610 546854
rect 219846 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 250330 546854
rect 250566 546618 281050 546854
rect 281286 546618 311770 546854
rect 312006 546618 342490 546854
rect 342726 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 373210 546854
rect 373446 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 420328 546854
rect 420564 546618 556056 546854
rect 556292 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 21008 543454
rect 21244 543218 155376 543454
rect 155612 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 204250 543454
rect 204486 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 234970 543454
rect 235206 543218 265690 543454
rect 265926 543218 296410 543454
rect 296646 543218 327130 543454
rect 327366 543218 357850 543454
rect 358086 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 421008 543454
rect 421244 543218 555376 543454
rect 555612 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 21008 543134
rect 21244 542898 155376 543134
rect 155612 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 204250 543134
rect 204486 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 234970 543134
rect 235206 542898 265690 543134
rect 265926 542898 296410 543134
rect 296646 542898 327130 543134
rect 327366 542898 357850 543134
rect 358086 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 421008 543134
rect 421244 542898 555376 543134
rect 555612 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 20328 511174
rect 20564 510938 156056 511174
rect 156292 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 219610 511174
rect 219846 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 250330 511174
rect 250566 510938 281050 511174
rect 281286 510938 311770 511174
rect 312006 510938 342490 511174
rect 342726 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 373210 511174
rect 373446 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 420328 511174
rect 420564 510938 556056 511174
rect 556292 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 20328 510854
rect 20564 510618 156056 510854
rect 156292 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 219610 510854
rect 219846 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 250330 510854
rect 250566 510618 281050 510854
rect 281286 510618 311770 510854
rect 312006 510618 342490 510854
rect 342726 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 373210 510854
rect 373446 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 420328 510854
rect 420564 510618 556056 510854
rect 556292 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 21008 507454
rect 21244 507218 155376 507454
rect 155612 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 204250 507454
rect 204486 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 234970 507454
rect 235206 507218 265690 507454
rect 265926 507218 296410 507454
rect 296646 507218 327130 507454
rect 327366 507218 357850 507454
rect 358086 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 421008 507454
rect 421244 507218 555376 507454
rect 555612 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 21008 507134
rect 21244 506898 155376 507134
rect 155612 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 204250 507134
rect 204486 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 234970 507134
rect 235206 506898 265690 507134
rect 265926 506898 296410 507134
rect 296646 506898 327130 507134
rect 327366 506898 357850 507134
rect 358086 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 421008 507134
rect 421244 506898 555376 507134
rect 555612 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 279866 497494
rect 280102 497258 280186 497494
rect 280422 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 279866 497174
rect 280102 496938 280186 497174
rect 280422 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 276146 493774
rect 276382 493538 276466 493774
rect 276702 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 276146 493454
rect 276382 493218 276466 493454
rect 276702 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 272426 490054
rect 272662 489818 272746 490054
rect 272982 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 272426 489734
rect 272662 489498 272746 489734
rect 272982 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 209610 439174
rect 209846 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 240330 439174
rect 240566 438938 271050 439174
rect 271286 438938 301770 439174
rect 302006 438938 332490 439174
rect 332726 438938 363210 439174
rect 363446 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 209610 438854
rect 209846 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 240330 438854
rect 240566 438618 271050 438854
rect 271286 438618 301770 438854
rect 302006 438618 332490 438854
rect 332726 438618 363210 438854
rect 363446 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 194250 435454
rect 194486 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 224970 435454
rect 225206 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 255690 435454
rect 255926 435218 286410 435454
rect 286646 435218 317130 435454
rect 317366 435218 347850 435454
rect 348086 435218 378570 435454
rect 378806 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 194250 435134
rect 194486 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 224970 435134
rect 225206 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 255690 435134
rect 255926 434898 286410 435134
rect 286646 434898 317130 435134
rect 317366 434898 347850 435134
rect 348086 434898 378570 435134
rect 378806 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 209610 403174
rect 209846 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 240330 403174
rect 240566 402938 271050 403174
rect 271286 402938 301770 403174
rect 302006 402938 332490 403174
rect 332726 402938 363210 403174
rect 363446 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 209610 402854
rect 209846 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 240330 402854
rect 240566 402618 271050 402854
rect 271286 402618 301770 402854
rect 302006 402618 332490 402854
rect 332726 402618 363210 402854
rect 363446 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 194250 399454
rect 194486 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 224970 399454
rect 225206 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 255690 399454
rect 255926 399218 286410 399454
rect 286646 399218 317130 399454
rect 317366 399218 347850 399454
rect 348086 399218 378570 399454
rect 378806 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 194250 399134
rect 194486 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 224970 399134
rect 225206 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 255690 399134
rect 255926 398898 286410 399134
rect 286646 398898 317130 399134
rect 317366 398898 347850 399134
rect 348086 398898 378570 399134
rect 378806 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 209610 367174
rect 209846 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 240330 367174
rect 240566 366938 271050 367174
rect 271286 366938 301770 367174
rect 302006 366938 332490 367174
rect 332726 366938 363210 367174
rect 363446 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 209610 366854
rect 209846 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 240330 366854
rect 240566 366618 271050 366854
rect 271286 366618 301770 366854
rect 302006 366618 332490 366854
rect 332726 366618 363210 366854
rect 363446 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 194250 363454
rect 194486 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 224970 363454
rect 225206 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 255690 363454
rect 255926 363218 286410 363454
rect 286646 363218 317130 363454
rect 317366 363218 347850 363454
rect 348086 363218 378570 363454
rect 378806 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 194250 363134
rect 194486 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 224970 363134
rect 225206 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 255690 363134
rect 255926 362898 286410 363134
rect 286646 362898 317130 363134
rect 317366 362898 347850 363134
rect 348086 362898 378570 363134
rect 378806 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 209610 331174
rect 209846 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 240330 331174
rect 240566 330938 271050 331174
rect 271286 330938 301770 331174
rect 302006 330938 332490 331174
rect 332726 330938 363210 331174
rect 363446 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 209610 330854
rect 209846 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 240330 330854
rect 240566 330618 271050 330854
rect 271286 330618 301770 330854
rect 302006 330618 332490 330854
rect 332726 330618 363210 330854
rect 363446 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 194250 327454
rect 194486 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 224970 327454
rect 225206 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 255690 327454
rect 255926 327218 286410 327454
rect 286646 327218 317130 327454
rect 317366 327218 347850 327454
rect 348086 327218 378570 327454
rect 378806 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 194250 327134
rect 194486 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 224970 327134
rect 225206 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 255690 327134
rect 255926 326898 286410 327134
rect 286646 326898 317130 327134
rect 317366 326898 347850 327134
rect 348086 326898 378570 327134
rect 378806 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 209610 295174
rect 209846 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 240330 295174
rect 240566 294938 271050 295174
rect 271286 294938 301770 295174
rect 302006 294938 332490 295174
rect 332726 294938 363210 295174
rect 363446 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 209610 294854
rect 209846 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 240330 294854
rect 240566 294618 271050 294854
rect 271286 294618 301770 294854
rect 302006 294618 332490 294854
rect 332726 294618 363210 294854
rect 363446 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 194250 291454
rect 194486 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 224970 291454
rect 225206 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 255690 291454
rect 255926 291218 286410 291454
rect 286646 291218 317130 291454
rect 317366 291218 347850 291454
rect 348086 291218 378570 291454
rect 378806 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 194250 291134
rect 194486 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 224970 291134
rect 225206 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 255690 291134
rect 255926 290898 286410 291134
rect 286646 290898 317130 291134
rect 317366 290898 347850 291134
rect 348086 290898 378570 291134
rect 378806 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 63866 281494
rect 64102 281258 64186 281494
rect 64422 281258 99866 281494
rect 100102 281258 100186 281494
rect 100422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 63866 281174
rect 64102 280938 64186 281174
rect 64422 280938 99866 281174
rect 100102 280938 100186 281174
rect 100422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 209610 259174
rect 209846 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 240330 259174
rect 240566 258938 271050 259174
rect 271286 258938 301770 259174
rect 302006 258938 332490 259174
rect 332726 258938 363210 259174
rect 363446 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 209610 258854
rect 209846 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 240330 258854
rect 240566 258618 271050 258854
rect 271286 258618 301770 258854
rect 302006 258618 332490 258854
rect 332726 258618 363210 258854
rect 363446 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 194250 255454
rect 194486 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 224970 255454
rect 225206 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 255690 255454
rect 255926 255218 286410 255454
rect 286646 255218 317130 255454
rect 317366 255218 347850 255454
rect 348086 255218 378570 255454
rect 378806 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 194250 255134
rect 194486 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 224970 255134
rect 225206 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 255690 255134
rect 255926 254898 286410 255134
rect 286646 254898 317130 255134
rect 317366 254898 347850 255134
rect 348086 254898 378570 255134
rect 378806 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 276146 241774
rect 276382 241538 276466 241774
rect 276702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 276146 241454
rect 276382 241218 276466 241454
rect 276702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 20328 187174
rect 20564 186938 156056 187174
rect 156292 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 420328 187174
rect 420564 186938 556056 187174
rect 556292 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 20328 186854
rect 20564 186618 156056 186854
rect 156292 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 420328 186854
rect 420564 186618 556056 186854
rect 556292 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 21008 183454
rect 21244 183218 155376 183454
rect 155612 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 421008 183454
rect 421244 183218 555376 183454
rect 555612 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 21008 183134
rect 21244 182898 155376 183134
rect 155612 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 421008 183134
rect 421244 182898 555376 183134
rect 555612 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 20328 151174
rect 20564 150938 156056 151174
rect 156292 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 420328 151174
rect 420564 150938 556056 151174
rect 556292 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 20328 150854
rect 20564 150618 156056 150854
rect 156292 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 420328 150854
rect 420564 150618 556056 150854
rect 556292 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 21008 147454
rect 21244 147218 155376 147454
rect 155612 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 421008 147454
rect 421244 147218 555376 147454
rect 555612 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 21008 147134
rect 21244 146898 155376 147134
rect 155612 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 421008 147134
rect 421244 146898 555376 147134
rect 555612 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 20328 115174
rect 20564 114938 156056 115174
rect 156292 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 420328 115174
rect 420564 114938 556056 115174
rect 556292 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 20328 114854
rect 20564 114618 156056 114854
rect 156292 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 420328 114854
rect 420564 114618 556056 114854
rect 556292 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111337 181826 111454
rect 2382 111218 21008 111337
rect -8726 111134 21008 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 111101 21008 111134
rect 21244 111101 155376 111337
rect 155612 111218 181826 111337
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111337 577826 111454
rect 398382 111218 421008 111337
rect 155612 111134 421008 111218
rect 155612 111101 181826 111134
rect 2382 110898 181826 111101
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 111101 421008 111134
rect 421244 111101 555376 111337
rect 555612 111218 577826 111337
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect 555612 111134 592650 111218
rect 555612 111101 577826 111134
rect 398382 110898 577826 111101
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 20328 79174
rect 20564 78938 156056 79174
rect 156292 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 220328 79174
rect 220564 78938 356056 79174
rect 356292 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 420328 79174
rect 420564 78938 556056 79174
rect 556292 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 20328 78854
rect 20564 78618 156056 78854
rect 156292 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 220328 78854
rect 220564 78618 356056 78854
rect 356292 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 420328 78854
rect 420564 78618 556056 78854
rect 556292 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 21008 75454
rect 21244 75218 155376 75454
rect 155612 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 221008 75454
rect 221244 75218 355376 75454
rect 355612 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 421008 75454
rect 421244 75218 555376 75454
rect 555612 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 21008 75134
rect 21244 74898 155376 75134
rect 155612 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 221008 75134
rect 221244 74898 355376 75134
rect 355612 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 421008 75134
rect 421244 74898 555376 75134
rect 555612 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 20328 43174
rect 20564 42938 156056 43174
rect 156292 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 220328 43174
rect 220564 42938 356056 43174
rect 356292 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 420328 43174
rect 420564 42938 556056 43174
rect 556292 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 20328 42854
rect 20564 42618 156056 42854
rect 156292 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 220328 42854
rect 220564 42618 356056 42854
rect 356292 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 420328 42854
rect 420564 42618 556056 42854
rect 556292 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 21008 39454
rect 21244 39218 155376 39454
rect 155612 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 221008 39454
rect 221244 39218 355376 39454
rect 355612 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 421008 39454
rect 421244 39218 555376 39454
rect 555612 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 21008 39134
rect 21244 38898 155376 39134
rect 155612 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 221008 39134
rect 221244 38898 355376 39134
rect 355612 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 421008 39134
rect 421244 38898 555376 39134
rect 555612 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18023 592650 18098
rect -8726 18014 52706 18023
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17787 52706 18014
rect 52942 17787 53026 18023
rect 53262 17787 88706 18023
rect 88942 17787 89026 18023
rect 89262 17787 124706 18023
rect 124942 17787 125026 18023
rect 125262 18014 232706 18023
rect 125262 17787 160706 18014
rect 17262 17778 160706 17787
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17787 232706 18014
rect 232942 17787 233026 18023
rect 233262 17787 304706 18023
rect 304942 17787 305026 18023
rect 305262 17787 340706 18023
rect 340942 17787 341026 18023
rect 341262 18014 484706 18023
rect 341262 17787 376706 18014
rect 197262 17778 376706 17787
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17787 484706 18014
rect 484942 17787 485026 18023
rect 485262 17787 556706 18023
rect 556942 17787 557026 18023
rect 557262 18014 592650 18023
rect 557262 17787 589182 18014
rect 413262 17778 589182 17787
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use io_interface  IO_interface
timestamp 0
transform 1 0 190000 0 1 250000
box 1066 0 198850 200000
use sky130_sram_2kbyte_1rw1r_32x512_8  data_memory
timestamp 0
transform 1 0 220000 0 1 20000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory0
timestamp 0
transform 1 0 420000 0 1 110000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory1
timestamp 0
transform 1 0 420000 0 1 500000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory2
timestamp 0
transform 1 0 20000 0 1 110000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory3
timestamp 0
transform 1 0 20000 0 1 500000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory4
timestamp 0
transform 1 0 420000 0 1 20000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory5
timestamp 0
transform 1 0 420000 0 1 590000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory6
timestamp 0
transform 1 0 20000 0 1 20000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  instr_memory7
timestamp 0
transform 1 0 20000 0 1 590000
box 0 0 136620 83308
use processor  uP
timestamp 0
transform 1 0 200000 0 1 500000
box 1066 0 178886 180000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 17940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 195244 38414 497940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 675244 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 17940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 195244 74414 497940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 675244 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 18064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 195244 110414 498064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 675244 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 18064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 195244 146414 498064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 675244 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 18064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 105244 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 18064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 105244 254414 501375 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 678961 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 18064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 105244 290414 249743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 678961 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 17940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 105244 326414 249743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 678961 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 249743 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 451537 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 18064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 195244 434414 498064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 675244 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 17940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 195244 470414 497940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 675244 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 17940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 195244 506414 497940 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 675244 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 18064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 195244 542414 498064 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 675244 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 17940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 195244 45854 497940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 675244 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 18064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 195244 81854 498064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 675244 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 18064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 195244 117854 498064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 675244 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 18064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 195244 153854 498064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 675244 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 18064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 105244 225854 250068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 449580 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 17940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 105244 261854 249743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 678961 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 18064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 105244 297854 249743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 678961 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 18064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 105244 333854 249743 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 451537 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 17940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 195244 441854 497940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 675244 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 18064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 195244 477854 498064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 675244 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 17940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 195244 513854 497940 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 675244 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 18064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 195244 549854 498064 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 675244 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 18064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 195244 53294 498064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 18064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 195244 89294 498064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 18064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 195244 125294 498064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 18064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 105244 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 17940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 105244 269294 249743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 18064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 105244 305294 249743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 18064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 105244 341294 249743 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 451537 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 17940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 195244 449294 497940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 18064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 195244 485294 498064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 17940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 195244 521294 497940 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 18064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 195244 557294 498064 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 195244 24734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 195244 60734 497940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 195244 96734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 195244 132734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 105244 240734 250068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 449580 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 105244 276734 249743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 451537 276734 501375 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 105244 312734 249743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 451537 312734 501375 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 105244 348734 249743 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 451537 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 195244 420734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 195244 456734 497940 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 195244 492734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 195244 528734 498064 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 195244 21014 498064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 195244 57014 497940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 195244 93014 498064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 195244 129014 498064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 105244 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 105244 273014 249743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 451537 273014 501375 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 105244 309014 249743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 451537 309014 501375 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 105244 345014 249743 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 451537 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 195244 453014 497940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 195244 489014 497940 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 195244 525014 498064 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 195244 28454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 675244 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 195244 64454 497940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 675244 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 195244 100454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 675244 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 195244 136454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 675244 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 105244 244454 501375 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 105244 280454 249743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 451537 280454 501375 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 105244 316454 249743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 451537 316454 501375 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 105244 352454 249743 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 451537 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 195244 424454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 675244 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 195244 460454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 675244 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 195244 496454 497940 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 675244 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 195244 532454 498064 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 675244 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 17940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 195244 42134 497940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 675244 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 17940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 195244 78134 497940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 675244 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 17940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 195244 114134 497940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 675244 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 18064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 195244 150134 498064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 675244 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 18064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 105244 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 17940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 105244 258134 249743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 678961 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 17940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 105244 294134 249743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 678961 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 18064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 105244 330134 249743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 678961 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 249743 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 451537 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 18064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 195244 438134 498064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 675244 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 17940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 195244 474134 497940 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 675244 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 18064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 195244 510134 498064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 675244 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 18064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 195244 546134 498064 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 675244 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 18064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 195244 49574 498064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 675244 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 18064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 195244 85574 498064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 675244 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 17940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 195244 121574 497940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 675244 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 18064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 195244 157574 498064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 675244 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 18064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 105244 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 17940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 105244 265574 249743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 678961 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 17940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 105244 301574 249743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 678961 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 18064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 105244 337574 249743 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 451537 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 500068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 679452 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 17940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 195244 445574 497940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 675244 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 17940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 195244 481574 497940 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 675244 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 18064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 195244 517574 498064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 675244 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 18064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 195244 553574 498064 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 675244 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 155494 651336 155494 651336 0 vccd1
rlabel via4 369704 658776 369704 658776 0 vccd2
rlabel via4 377144 666216 377144 666216 0 vdda1
rlabel via4 348584 673656 348584 673656 0 vdda2
rlabel via4 344864 669936 344864 669936 0 vssa1
rlabel via4 352304 677376 352304 677376 0 vssa2
rlabel via4 156174 655056 156174 655056 0 vssd1
rlabel via4 337424 662496 337424 662496 0 vssd2
rlabel metal1 386492 248370 386492 248370 0 Serial_input
rlabel metal1 387228 248302 387228 248302 0 Serial_output
rlabel metal3 19719 118334 19719 118334 0 clk
rlabel metal2 236026 18513 236026 18513 0 data_mem_addr\[0\]
rlabel metal4 237084 19040 237084 19040 0 data_mem_addr\[1\]
rlabel via2 216706 48229 216706 48229 0 data_mem_addr\[2\]
rlabel metal2 216706 50507 216706 50507 0 data_mem_addr\[3\]
rlabel metal2 216798 51731 216798 51731 0 data_mem_addr\[4\]
rlabel via1 268594 449565 268594 449565 0 data_mem_addr\[5\]
rlabel metal2 269882 450218 269882 450218 0 data_mem_addr\[6\]
rlabel metal2 216706 56253 216706 56253 0 data_mem_addr\[7\]
rlabel metal3 217281 28492 217281 28492 0 data_mem_csb
rlabel metal1 188554 447950 188554 447950 0 data_read_data\[0\]
rlabel metal2 273286 17833 273286 17833 0 data_read_data\[10\]
rlabel metal4 276092 18292 276092 18292 0 data_read_data\[11\]
rlabel metal4 277196 18632 277196 18632 0 data_read_data\[12\]
rlabel metal2 275770 450864 275770 450864 0 data_read_data\[13\]
rlabel metal2 218730 133790 218730 133790 0 data_read_data\[14\]
rlabel metal2 277242 451068 277242 451068 0 data_read_data\[15\]
rlabel metal2 250654 18921 250654 18921 0 data_read_data\[1\]
rlabel metal2 253598 18785 253598 18785 0 data_read_data\[2\]
rlabel via2 255990 18683 255990 18683 0 data_read_data\[3\]
rlabel metal2 267897 449956 267897 449956 0 data_read_data\[4\]
rlabel metal2 269146 454944 269146 454944 0 data_read_data\[5\]
rlabel metal2 270105 449956 270105 449956 0 data_read_data\[6\]
rlabel metal2 271209 449956 271209 449956 0 data_read_data\[7\]
rlabel metal4 268364 18632 268364 18632 0 data_read_data\[8\]
rlabel via2 270526 17595 270526 17595 0 data_read_data\[9\]
rlabel metal4 238188 19108 238188 19108 0 data_wmask\[0\]
rlabel metal4 239660 19380 239660 19380 0 data_wmask\[1\]
rlabel metal4 240580 19448 240580 19448 0 data_wmask\[2\]
rlabel metal4 241684 19312 241684 19312 0 data_wmask\[3\]
rlabel via2 243110 18547 243110 18547 0 data_write_data\[0\]
rlabel metal4 254564 18632 254564 18632 0 data_write_data\[10\]
rlabel metal2 255346 17255 255346 17255 0 data_write_data\[11\]
rlabel metal2 256726 17289 256726 17289 0 data_write_data\[12\]
rlabel metal2 276191 449956 276191 449956 0 data_write_data\[13\]
rlabel metal2 276729 449956 276729 449956 0 data_write_data\[14\]
rlabel metal2 259578 17527 259578 17527 0 data_write_data\[15\]
rlabel via2 244306 19261 244306 19261 0 data_write_data\[1\]
rlabel metal2 245318 19193 245318 19193 0 data_write_data\[2\]
rlabel via2 246422 19227 246422 19227 0 data_write_data\[3\]
rlabel metal2 268265 449956 268265 449956 0 data_write_data\[4\]
rlabel metal4 248676 18496 248676 18496 0 data_write_data\[5\]
rlabel metal2 250102 19057 250102 19057 0 data_write_data\[6\]
rlabel via2 251206 17051 251206 17051 0 data_write_data\[7\]
rlabel via2 252310 18819 252310 18819 0 data_write_data\[8\]
rlabel metal3 191797 369852 191797 369852 0 data_write_data\[9\]
rlabel metal2 277833 449956 277833 449956 0 dataw_enb
rlabel metal2 372462 680959 372462 680959 0 hlt
rlabel metal4 35972 18292 35972 18292 0 instr_mem_addr_9bit\[0\]
rlabel via2 36570 17901 36570 17901 0 instr_mem_addr_9bit\[1\]
rlabel via2 17894 138261 17894 138261 0 instr_mem_addr_9bit\[2\]
rlabel metal3 19719 139958 19719 139958 0 instr_mem_addr_9bit\[3\]
rlabel metal3 17342 140828 17342 140828 0 instr_mem_addr_9bit\[4\]
rlabel metal3 19719 622814 19719 622814 0 instr_mem_addr_9bit\[5\]
rlabel metal3 19719 623766 19719 623766 0 instr_mem_addr_9bit\[6\]
rlabel metal3 19719 55942 19719 55942 0 instr_mem_addr_9bit\[7\]
rlabel metal3 19719 56894 19719 56894 0 instr_mem_addr_9bit\[8\]
rlabel metal2 308522 451136 308522 451136 0 instr_mem_csb\[0\]
rlabel metal2 304329 449956 304329 449956 0 instr_mem_csb\[1\]
rlabel metal3 19719 118062 19719 118062 0 instr_mem_csb\[2\]
rlabel metal3 19742 508062 19742 508062 0 instr_mem_csb\[3\]
rlabel metal2 291962 451442 291962 451442 0 instr_mem_csb\[4\]
rlabel metal2 287401 449956 287401 449956 0 instr_mem_csb\[5\]
rlabel metal3 19903 28062 19903 28062 0 instr_mem_csb\[6\]
rlabel metal3 19719 598062 19719 598062 0 instr_mem_csb\[7\]
rlabel metal2 390126 279905 390126 279905 0 instr_read_data0\[0\]
rlabel metal2 319194 450847 319194 450847 0 instr_read_data0\[10\]
rlabel metal2 388838 280432 388838 280432 0 instr_read_data0\[11\]
rlabel metal2 418830 280109 418830 280109 0 instr_read_data0\[12\]
rlabel metal4 480966 109948 480966 109948 0 instr_read_data0\[13\]
rlabel metal2 332442 450048 332442 450048 0 instr_read_data0\[14\]
rlabel metal4 485998 109948 485998 109948 0 instr_read_data0\[15\]
rlabel metal4 488310 109948 488310 109948 0 instr_read_data0\[16\]
rlabel metal2 342010 450422 342010 450422 0 instr_read_data0\[17\]
rlabel metal2 344954 451578 344954 451578 0 instr_read_data0\[18\]
rlabel metal2 347898 450116 347898 450116 0 instr_read_data0\[19\]
rlabel metal2 392610 280194 392610 280194 0 instr_read_data0\[1\]
rlabel metal2 350842 450150 350842 450150 0 instr_read_data0\[20\]
rlabel metal2 353786 450184 353786 450184 0 instr_read_data0\[21\]
rlabel metal4 503542 109948 503542 109948 0 instr_read_data0\[22\]
rlabel metal2 410826 279616 410826 279616 0 instr_read_data0\[23\]
rlabel metal2 410734 281214 410734 281214 0 instr_read_data0\[24\]
rlabel via1 365746 449939 365746 449939 0 instr_read_data0\[25\]
rlabel metal2 368506 450286 368506 450286 0 instr_read_data0\[26\]
rlabel metal2 411010 279582 411010 279582 0 instr_read_data0\[27\]
rlabel metal2 411102 279582 411102 279582 0 instr_read_data0\[28\]
rlabel metal4 520950 109948 520950 109948 0 instr_read_data0\[29\]
rlabel metal2 287914 450643 287914 450643 0 instr_read_data0\[2\]
rlabel metal2 388654 280092 388654 280092 0 instr_read_data0\[30\]
rlabel metal4 525982 109948 525982 109948 0 instr_read_data0\[31\]
rlabel metal2 292330 450779 292330 450779 0 instr_read_data0\[3\]
rlabel metal2 408158 279089 408158 279089 0 instr_read_data0\[4\]
rlabel metal2 408342 280024 408342 280024 0 instr_read_data0\[5\]
rlabel metal2 388746 278664 388746 278664 0 instr_read_data0\[6\]
rlabel via1 309074 449565 309074 449565 0 instr_read_data0\[7\]
rlabel via1 312846 449667 312846 449667 0 instr_read_data0\[8\]
rlabel metal2 315882 451510 315882 451510 0 instr_read_data0\[9\]
rlabel metal4 448326 499818 448326 499818 0 instr_read_data1\[0\]
rlabel metal2 319417 449956 319417 449956 0 instr_read_data1\[10\]
rlabel metal1 398866 476782 398866 476782 0 instr_read_data1\[11\]
rlabel metal4 478518 499818 478518 499818 0 instr_read_data1\[12\]
rlabel metal4 480966 499818 480966 499818 0 instr_read_data1\[13\]
rlabel metal2 332757 449956 332757 449956 0 instr_read_data1\[14\]
rlabel metal4 485998 499818 485998 499818 0 instr_read_data1\[15\]
rlabel metal4 488310 499818 488310 499818 0 instr_read_data1\[16\]
rlabel metal2 342325 449956 342325 449956 0 instr_read_data1\[17\]
rlabel metal2 345177 449956 345177 449956 0 instr_read_data1\[18\]
rlabel metal2 348121 449956 348121 449956 0 instr_read_data1\[19\]
rlabel metal4 450774 499818 450774 499818 0 instr_read_data1\[1\]
rlabel metal2 351065 449956 351065 449956 0 instr_read_data1\[20\]
rlabel metal2 354009 449956 354009 449956 0 instr_read_data1\[21\]
rlabel metal4 503542 499818 503542 499818 0 instr_read_data1\[22\]
rlabel metal4 505990 499818 505990 499818 0 instr_read_data1\[23\]
rlabel metal4 508574 499818 508574 499818 0 instr_read_data1\[24\]
rlabel metal2 365930 457868 365930 457868 0 instr_read_data1\[25\]
rlabel metal2 368729 449956 368729 449956 0 instr_read_data1\[26\]
rlabel metal2 371358 465383 371358 465383 0 instr_read_data1\[27\]
rlabel metal1 445786 464406 445786 464406 0 instr_read_data1\[28\]
rlabel metal4 520950 499818 520950 499818 0 instr_read_data1\[29\]
rlabel metal2 288137 449956 288137 449956 0 instr_read_data1\[2\]
rlabel metal4 523398 499818 523398 499818 0 instr_read_data1\[30\]
rlabel metal4 525982 499818 525982 499818 0 instr_read_data1\[31\]
rlabel metal1 374210 488002 374210 488002 0 instr_read_data1\[3\]
rlabel metal1 377568 483786 377568 483786 0 instr_read_data1\[4\]
rlabel metal4 461110 499818 461110 499818 0 instr_read_data1\[5\]
rlabel metal4 463558 499818 463558 499818 0 instr_read_data1\[6\]
rlabel metal2 309205 449956 309205 449956 0 instr_read_data1\[7\]
rlabel metal2 312793 449956 312793 449956 0 instr_read_data1\[8\]
rlabel metal2 316151 449956 316151 449956 0 instr_read_data1\[9\]
rlabel metal2 279673 449956 279673 449956 0 instr_read_data2\[0\]
rlabel metal2 319785 449956 319785 449956 0 instr_read_data2\[10\]
rlabel metal4 76070 109948 76070 109948 0 instr_read_data2\[11\]
rlabel metal4 78518 109948 78518 109948 0 instr_read_data2\[12\]
rlabel metal4 80966 109948 80966 109948 0 instr_read_data2\[13\]
rlabel metal2 333033 449956 333033 449956 0 instr_read_data2\[14\]
rlabel metal2 158194 278664 158194 278664 0 instr_read_data2\[15\]
rlabel metal2 156630 279072 156630 279072 0 instr_read_data2\[16\]
rlabel metal2 342647 449956 342647 449956 0 instr_read_data2\[17\]
rlabel metal2 345690 450456 345690 450456 0 instr_read_data2\[18\]
rlabel metal2 348489 449956 348489 449956 0 instr_read_data2\[19\]
rlabel metal4 50774 109812 50774 109812 0 instr_read_data2\[1\]
rlabel metal2 351578 450388 351578 450388 0 instr_read_data2\[20\]
rlabel metal2 354522 450031 354522 450031 0 instr_read_data2\[21\]
rlabel metal3 192901 450500 192901 450500 0 instr_read_data2\[22\]
rlabel metal2 360311 449956 360311 449956 0 instr_read_data2\[23\]
rlabel metal2 363255 449956 363255 449956 0 instr_read_data2\[24\]
rlabel metal2 366153 449956 366153 449956 0 instr_read_data2\[25\]
rlabel metal2 369097 449956 369097 449956 0 instr_read_data2\[26\]
rlabel metal4 115918 109948 115918 109948 0 instr_read_data2\[27\]
rlabel metal4 118502 109948 118502 109948 0 instr_read_data2\[28\]
rlabel metal4 120950 109948 120950 109948 0 instr_read_data2\[29\]
rlabel metal2 288650 450150 288650 450150 0 instr_read_data2\[2\]
rlabel metal2 381071 449956 381071 449956 0 instr_read_data2\[30\]
rlabel metal3 386607 449684 386607 449684 0 instr_read_data2\[31\]
rlabel metal4 56078 109812 56078 109812 0 instr_read_data2\[3\]
rlabel metal4 58526 109948 58526 109948 0 instr_read_data2\[4\]
rlabel metal4 61110 109812 61110 109812 0 instr_read_data2\[5\]
rlabel metal4 63558 109948 63558 109948 0 instr_read_data2\[6\]
rlabel metal2 309481 449956 309481 449956 0 instr_read_data2\[7\]
rlabel metal2 313214 458303 313214 458303 0 instr_read_data2\[8\]
rlabel metal3 192901 450772 192901 450772 0 instr_read_data2\[9\]
rlabel metal2 280239 449956 280239 449956 0 instr_read_data3\[0\]
rlabel metal4 73622 499818 73622 499818 0 instr_read_data3\[10\]
rlabel metal4 76070 499818 76070 499818 0 instr_read_data3\[11\]
rlabel metal4 78518 499818 78518 499818 0 instr_read_data3\[12\]
rlabel metal4 80966 499818 80966 499818 0 instr_read_data3\[13\]
rlabel metal2 333401 449956 333401 449956 0 instr_read_data3\[14\]
rlabel metal1 211876 483718 211876 483718 0 instr_read_data3\[15\]
rlabel metal2 340025 449956 340025 449956 0 instr_read_data3\[16\]
rlabel metal2 342969 449956 342969 449956 0 instr_read_data3\[17\]
rlabel metal2 345913 449956 345913 449956 0 instr_read_data3\[18\]
rlabel metal2 348857 449956 348857 449956 0 instr_read_data3\[19\]
rlabel metal4 50774 499818 50774 499818 0 instr_read_data3\[1\]
rlabel metal2 351999 449956 351999 449956 0 instr_read_data3\[20\]
rlabel metal4 100958 499818 100958 499818 0 instr_read_data3\[21\]
rlabel metal4 103316 498168 103316 498168 0 instr_read_data3\[22\]
rlabel metal2 360633 449956 360633 449956 0 instr_read_data3\[23\]
rlabel metal2 363577 449956 363577 449956 0 instr_read_data3\[24\]
rlabel metal2 366521 449956 366521 449956 0 instr_read_data3\[25\]
rlabel metal2 369465 449956 369465 449956 0 instr_read_data3\[26\]
rlabel metal4 115918 499818 115918 499818 0 instr_read_data3\[27\]
rlabel metal4 118502 499818 118502 499818 0 instr_read_data3\[28\]
rlabel metal4 120950 499818 120950 499818 0 instr_read_data3\[29\]
rlabel metal2 288873 449956 288873 449956 0 instr_read_data3\[2\]
rlabel metal2 381287 449956 381287 449956 0 instr_read_data3\[30\]
rlabel metal2 384185 449956 384185 449956 0 instr_read_data3\[31\]
rlabel metal4 56078 499818 56078 499818 0 instr_read_data3\[3\]
rlabel metal4 58526 499818 58526 499818 0 instr_read_data3\[4\]
rlabel metal4 61110 499818 61110 499818 0 instr_read_data3\[5\]
rlabel metal4 63558 499818 63558 499818 0 instr_read_data3\[6\]
rlabel metal2 309849 449956 309849 449956 0 instr_read_data3\[7\]
rlabel metal2 313529 449956 313529 449956 0 instr_read_data3\[8\]
rlabel metal2 316841 449956 316841 449956 0 instr_read_data3\[9\]
rlabel metal2 447166 17459 447166 17459 0 instr_read_data4\[0\]
rlabel metal2 388470 234124 388470 234124 0 instr_read_data4\[10\]
rlabel metal2 407974 235705 407974 235705 0 instr_read_data4\[11\]
rlabel metal2 407790 235807 407790 235807 0 instr_read_data4\[12\]
rlabel metal4 480700 18564 480700 18564 0 instr_read_data4\[13\]
rlabel metal2 333769 449956 333769 449956 0 instr_read_data4\[14\]
rlabel metal4 485998 19773 485998 19773 0 instr_read_data4\[15\]
rlabel metal2 488290 19737 488290 19737 0 instr_read_data4\[16\]
rlabel metal2 405122 237184 405122 237184 0 instr_read_data4\[17\]
rlabel metal2 346426 451646 346426 451646 0 instr_read_data4\[18\]
rlabel via1 349646 449701 349646 449701 0 instr_read_data4\[19\]
rlabel metal2 449926 17391 449926 17391 0 instr_read_data4\[1\]
rlabel metal2 352314 450983 352314 450983 0 instr_read_data4\[20\]
rlabel metal2 500986 19465 500986 19465 0 instr_read_data4\[21\]
rlabel metal2 503562 19431 503562 19431 0 instr_read_data4\[22\]
rlabel via2 505862 18853 505862 18853 0 instr_read_data4\[23\]
rlabel via2 508438 18819 508438 18819 0 instr_read_data4\[24\]
rlabel metal4 511060 18020 511060 18020 0 instr_read_data4\[25\]
rlabel metal4 513452 19176 513452 19176 0 instr_read_data4\[26\]
rlabel via2 515798 18955 515798 18955 0 instr_read_data4\[27\]
rlabel metal4 518420 19244 518420 19244 0 instr_read_data4\[28\]
rlabel metal2 485070 19040 485070 19040 0 instr_read_data4\[29\]
rlabel metal2 289241 449956 289241 449956 0 instr_read_data4\[2\]
rlabel via2 523342 18683 523342 18683 0 instr_read_data4\[30\]
rlabel metal2 525918 18649 525918 18649 0 instr_read_data4\[31\]
rlabel metal2 410550 235960 410550 235960 0 instr_read_data4\[3\]
rlabel metal2 458390 17969 458390 17969 0 instr_read_data4\[4\]
rlabel metal4 461110 19773 461110 19773 0 instr_read_data4\[5\]
rlabel metal4 463588 19108 463588 19108 0 instr_read_data4\[6\]
rlabel metal2 310217 449956 310217 449956 0 instr_read_data4\[7\]
rlabel metal2 313897 449956 313897 449956 0 instr_read_data4\[8\]
rlabel metal2 317209 449956 317209 449956 0 instr_read_data4\[9\]
rlabel metal4 448326 589988 448326 589988 0 instr_read_data5\[0\]
rlabel metal2 320889 449956 320889 449956 0 instr_read_data5\[10\]
rlabel metal2 418738 543847 418738 543847 0 instr_read_data5\[11\]
rlabel metal2 419014 543813 419014 543813 0 instr_read_data5\[12\]
rlabel metal4 480966 589988 480966 589988 0 instr_read_data5\[13\]
rlabel metal2 334137 449956 334137 449956 0 instr_read_data5\[14\]
rlabel metal4 485998 589988 485998 589988 0 instr_read_data5\[15\]
rlabel metal4 488310 589988 488310 589988 0 instr_read_data5\[16\]
rlabel metal4 489716 587880 489716 587880 0 instr_read_data5\[17\]
rlabel metal2 346649 449956 346649 449956 0 instr_read_data5\[18\]
rlabel metal2 349593 449956 349593 449956 0 instr_read_data5\[19\]
rlabel metal4 450774 589988 450774 589988 0 instr_read_data5\[1\]
rlabel metal2 352537 449956 352537 449956 0 instr_read_data5\[20\]
rlabel metal4 500958 589988 500958 589988 0 instr_read_data5\[21\]
rlabel metal4 503542 589988 503542 589988 0 instr_read_data5\[22\]
rlabel metal4 505990 589988 505990 589988 0 instr_read_data5\[23\]
rlabel metal2 364458 451102 364458 451102 0 instr_read_data5\[24\]
rlabel metal2 367402 450966 367402 450966 0 instr_read_data5\[25\]
rlabel metal1 446200 585922 446200 585922 0 instr_read_data5\[26\]
rlabel metal3 444659 584324 444659 584324 0 instr_read_data5\[27\]
rlabel metal3 446936 585684 446936 585684 0 instr_read_data5\[28\]
rlabel metal4 520950 589988 520950 589988 0 instr_read_data5\[29\]
rlabel metal2 289609 449956 289609 449956 0 instr_read_data5\[2\]
rlabel metal4 523398 589988 523398 589988 0 instr_read_data5\[30\]
rlabel metal2 385066 517912 385066 517912 0 instr_read_data5\[31\]
rlabel metal1 354384 474130 354384 474130 0 instr_read_data5\[3\]
rlabel metal2 380190 524110 380190 524110 0 instr_read_data5\[4\]
rlabel metal4 461110 589988 461110 589988 0 instr_read_data5\[5\]
rlabel metal2 306682 451000 306682 451000 0 instr_read_data5\[6\]
rlabel metal2 310730 451034 310730 451034 0 instr_read_data5\[7\]
rlabel metal2 314265 449956 314265 449956 0 instr_read_data5\[8\]
rlabel metal4 470396 588200 470396 588200 0 instr_read_data5\[9\]
rlabel metal4 48300 18564 48300 18564 0 instr_read_data6\[0\]
rlabel via2 73738 18819 73738 18819 0 instr_read_data6\[10\]
rlabel metal2 76130 18921 76130 18921 0 instr_read_data6\[11\]
rlabel metal2 78614 17765 78614 17765 0 instr_read_data6\[12\]
rlabel via2 81098 18955 81098 18955 0 instr_read_data6\[13\]
rlabel metal2 83858 17561 83858 17561 0 instr_read_data6\[14\]
rlabel metal2 179170 239513 179170 239513 0 instr_read_data6\[15\]
rlabel metal2 178894 237898 178894 237898 0 instr_read_data6\[16\]
rlabel metal2 178618 239479 178618 239479 0 instr_read_data6\[17\]
rlabel metal2 347017 449956 347017 449956 0 instr_read_data6\[18\]
rlabel metal2 96002 19193 96002 19193 0 instr_read_data6\[19\]
rlabel metal2 176410 238085 176410 238085 0 instr_read_data6\[1\]
rlabel via2 99314 17323 99314 17323 0 instr_read_data6\[20\]
rlabel via2 100970 19227 100970 19227 0 instr_read_data6\[21\]
rlabel metal2 176226 239445 176226 239445 0 instr_read_data6\[22\]
rlabel metal2 176502 238527 176502 238527 0 instr_read_data6\[23\]
rlabel metal2 364681 449956 364681 449956 0 instr_read_data6\[24\]
rlabel metal2 367625 449956 367625 449956 0 instr_read_data6\[25\]
rlabel via2 113482 18411 113482 18411 0 instr_read_data6\[26\]
rlabel metal4 115828 18496 115828 18496 0 instr_read_data6\[27\]
rlabel metal4 118588 19312 118588 19312 0 instr_read_data6\[28\]
rlabel metal4 120980 19244 120980 19244 0 instr_read_data6\[29\]
rlabel metal2 290069 449956 290069 449956 0 instr_read_data6\[2\]
rlabel metal4 122636 18428 122636 18428 0 instr_read_data6\[30\]
rlabel metal1 386768 451282 386768 451282 0 instr_read_data6\[31\]
rlabel metal2 56074 18785 56074 18785 0 instr_read_data6\[3\]
rlabel metal4 58604 18224 58604 18224 0 instr_read_data6\[4\]
rlabel via2 62054 17901 62054 17901 0 instr_read_data6\[5\]
rlabel via2 64722 17867 64722 17867 0 instr_read_data6\[6\]
rlabel metal2 310953 449956 310953 449956 0 instr_read_data6\[7\]
rlabel metal2 314778 450031 314778 450031 0 instr_read_data6\[8\]
rlabel via2 71714 17187 71714 17187 0 instr_read_data6\[9\]
rlabel metal1 241132 463318 241132 463318 0 instr_read_data7\[0\]
rlabel metal2 158010 526966 158010 526966 0 instr_read_data7\[10\]
rlabel metal4 76070 589852 76070 589852 0 instr_read_data7\[11\]
rlabel metal4 78518 589852 78518 589852 0 instr_read_data7\[12\]
rlabel metal2 331607 449956 331607 449956 0 instr_read_data7\[13\]
rlabel metal2 334873 449956 334873 449956 0 instr_read_data7\[14\]
rlabel metal4 195132 531352 195132 531352 0 instr_read_data7\[15\]
rlabel metal2 159390 533256 159390 533256 0 instr_read_data7\[16\]
rlabel metal2 344441 449956 344441 449956 0 instr_read_data7\[17\]
rlabel metal2 347385 449956 347385 449956 0 instr_read_data7\[18\]
rlabel metal2 350329 449956 350329 449956 0 instr_read_data7\[19\]
rlabel metal2 286074 450184 286074 450184 0 instr_read_data7\[1\]
rlabel metal4 98510 589988 98510 589988 0 instr_read_data7\[20\]
rlabel metal4 100958 589988 100958 589988 0 instr_read_data7\[21\]
rlabel metal4 103316 588880 103316 588880 0 instr_read_data7\[22\]
rlabel metal1 153272 585038 153272 585038 0 instr_read_data7\[23\]
rlabel metal2 365049 449956 365049 449956 0 instr_read_data7\[24\]
rlabel metal2 367993 449956 367993 449956 0 instr_read_data7\[25\]
rlabel metal4 113470 589988 113470 589988 0 instr_read_data7\[26\]
rlabel metal4 115918 589988 115918 589988 0 instr_read_data7\[27\]
rlabel metal4 199916 523600 199916 523600 0 instr_read_data7\[28\]
rlabel metal4 120950 589988 120950 589988 0 instr_read_data7\[29\]
rlabel metal2 290345 449956 290345 449956 0 instr_read_data7\[2\]
rlabel metal4 122636 588220 122636 588220 0 instr_read_data7\[30\]
rlabel metal2 385657 449956 385657 449956 0 instr_read_data7\[31\]
rlabel metal4 56078 589668 56078 589668 0 instr_read_data7\[3\]
rlabel metal4 58526 589988 58526 589988 0 instr_read_data7\[4\]
rlabel metal2 303225 449956 303225 449956 0 instr_read_data7\[5\]
rlabel metal2 307273 449956 307273 449956 0 instr_read_data7\[6\]
rlabel metal2 311321 449956 311321 449956 0 instr_read_data7\[7\]
rlabel metal2 315047 449956 315047 449956 0 instr_read_data7\[8\]
rlabel metal2 318313 449956 318313 449956 0 instr_read_data7\[9\]
rlabel metal4 38548 18428 38548 18428 0 instr_wmask\[0\]
rlabel metal2 38686 17153 38686 17153 0 instr_wmask\[1\]
rlabel metal4 40572 18496 40572 18496 0 instr_wmask\[2\]
rlabel metal3 41676 17952 41676 17952 0 instr_wmask\[3\]
rlabel metal1 41446 17102 41446 17102 0 instr_write_data\[0\]
rlabel metal2 18630 61710 18630 61710 0 instr_write_data\[10\]
rlabel metal2 56534 17306 56534 17306 0 instr_write_data\[11\]
rlabel metal2 57914 17051 57914 17051 0 instr_write_data\[12\]
rlabel metal4 58118 19705 58118 19705 0 instr_write_data\[13\]
rlabel metal4 59478 19705 59478 19705 0 instr_write_data\[14\]
rlabel metal4 60702 19705 60702 19705 0 instr_write_data\[15\]
rlabel metal1 41906 17170 41906 17170 0 instr_write_data\[1\]
rlabel metal1 42274 17238 42274 17238 0 instr_write_data\[2\]
rlabel metal4 446558 19705 446558 19705 0 instr_write_data\[3\]
rlabel metal4 447646 19841 447646 19841 0 instr_write_data\[4\]
rlabel metal4 448734 19841 448734 19841 0 instr_write_data\[5\]
rlabel metal2 307931 449956 307931 449956 0 instr_write_data\[6\]
rlabel metal1 20194 499970 20194 499970 0 instr_write_data\[7\]
rlabel metal2 315369 449956 315369 449956 0 instr_write_data\[8\]
rlabel metal4 53494 19773 53494 19773 0 instr_write_data\[9\]
rlabel metal3 19719 119966 19719 119966 0 instrw_enb
rlabel metal3 581908 6596 581908 6596 0 io_in[0]
rlabel metal2 580198 457079 580198 457079 0 io_in[10]
rlabel metal2 558302 492320 558302 492320 0 io_in[11]
rlabel metal2 579830 563703 579830 563703 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel metal2 565110 564128 565110 564128 0 io_in[14]
rlabel metal2 210167 449956 210167 449956 0 io_in[15]
rlabel metal2 211271 449956 211271 449956 0 io_in[16]
rlabel metal2 212329 449956 212329 449956 0 io_in[17]
rlabel metal2 213433 449956 213433 449956 0 io_in[18]
rlabel metal2 214537 449956 214537 449956 0 io_in[19]
rlabel metal2 194711 449956 194711 449956 0 io_in[1]
rlabel metal2 215641 449956 215641 449956 0 io_in[20]
rlabel metal2 216890 455896 216890 455896 0 io_in[21]
rlabel metal2 217849 449956 217849 449956 0 io_in[22]
rlabel metal2 218953 449956 218953 449956 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal3 1556 632060 1556 632060 0 io_in[25]
rlabel metal3 1832 579972 1832 579972 0 io_in[26]
rlabel metal3 1648 527884 1648 527884 0 io_in[27]
rlabel metal3 1694 475660 1694 475660 0 io_in[28]
rlabel metal3 475 423572 475 423572 0 io_in[29]
rlabel metal3 193775 451316 193775 451316 0 io_in[2]
rlabel metal3 1694 371348 1694 371348 0 io_in[30]
rlabel metal3 1648 319260 1648 319260 0 io_in[31]
rlabel metal3 1786 267172 1786 267172 0 io_in[32]
rlabel metal3 1832 214948 1832 214948 0 io_in[33]
rlabel metal3 1970 162860 1970 162860 0 io_in[34]
rlabel metal3 1832 110636 1832 110636 0 io_in[35]
rlabel metal3 1832 71604 1832 71604 0 io_in[36]
rlabel metal3 1832 32436 1832 32436 0 io_in[37]
rlabel metal2 566490 290479 566490 290479 0 io_in[3]
rlabel metal2 580198 166413 580198 166413 0 io_in[4]
rlabel metal2 579830 206329 579830 206329 0 io_in[5]
rlabel metal2 392702 350030 392702 350030 0 io_in[6]
rlabel metal2 390402 437189 390402 437189 0 io_in[7]
rlabel metal2 580198 352563 580198 352563 0 io_in[8]
rlabel metal1 388378 449786 388378 449786 0 io_in[9]
rlabel via3 194051 449276 194051 449276 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 566490 509558 566490 509558 0 io_oeb[11]
rlabel metal2 558210 544782 558210 544782 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 210489 449956 210489 449956 0 io_oeb[15]
rlabel metal2 211593 449956 211593 449956 0 io_oeb[16]
rlabel metal2 212789 449956 212789 449956 0 io_oeb[17]
rlabel metal2 332534 702093 332534 702093 0 io_oeb[18]
rlabel metal2 214905 449956 214905 449956 0 io_oeb[19]
rlabel metal2 195178 450711 195178 450711 0 io_oeb[1]
rlabel metal2 216009 449956 216009 449956 0 io_oeb[20]
rlabel metal2 217113 449956 217113 449956 0 io_oeb[21]
rlabel metal2 218217 449956 218217 449956 0 io_oeb[22]
rlabel metal1 11316 700230 11316 700230 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 1786 606084 1786 606084 0 io_oeb[25]
rlabel metal3 1832 553860 1832 553860 0 io_oeb[26]
rlabel metal3 1832 501772 1832 501772 0 io_oeb[27]
rlabel metal3 1832 449548 1832 449548 0 io_oeb[28]
rlabel metal3 1832 397460 1832 397460 0 io_oeb[29]
rlabel metal2 580014 112965 580014 112965 0 io_oeb[2]
rlabel metal3 1832 345372 1832 345372 0 io_oeb[30]
rlabel metal3 1602 293148 1602 293148 0 io_oeb[31]
rlabel metal3 1786 241060 1786 241060 0 io_oeb[32]
rlabel metal3 1832 188836 1832 188836 0 io_oeb[33]
rlabel metal3 1694 136748 1694 136748 0 io_oeb[34]
rlabel metal3 2016 84660 2016 84660 0 io_oeb[35]
rlabel metal3 1832 45492 1832 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal2 579646 192831 579646 192831 0 io_oeb[4]
rlabel metal3 582138 232356 582138 232356 0 io_oeb[5]
rlabel metal2 580198 272697 580198 272697 0 io_oeb[6]
rlabel metal2 391322 390660 391322 390660 0 io_oeb[7]
rlabel metal2 390310 417010 390310 417010 0 io_oeb[8]
rlabel metal3 582184 431596 582184 431596 0 io_oeb[9]
rlabel metal3 194005 450228 194005 450228 0 io_out[0]
rlabel metal2 580014 471019 580014 471019 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal2 580198 577269 580198 577269 0 io_out[12]
rlabel metal2 580198 630751 580198 630751 0 io_out[13]
rlabel metal2 209845 449956 209845 449956 0 io_out[14]
rlabel metal2 210857 449956 210857 449956 0 io_out[15]
rlabel metal2 211961 449956 211961 449956 0 io_out[16]
rlabel metal2 213065 449956 213065 449956 0 io_out[17]
rlabel metal2 214169 449956 214169 449956 0 io_out[18]
rlabel metal1 215602 500786 215602 500786 0 io_out[19]
rlabel metal3 582000 59636 582000 59636 0 io_out[1]
rlabel metal2 216377 449956 216377 449956 0 io_out[20]
rlabel metal2 217481 449956 217481 449956 0 io_out[21]
rlabel metal2 218585 449956 218585 449956 0 io_out[22]
rlabel metal2 24334 701974 24334 701974 0 io_out[23]
rlabel metal3 1924 671228 1924 671228 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 1878 566916 1878 566916 0 io_out[26]
rlabel metal2 3588 480240 3588 480240 0 io_out[27]
rlabel metal3 1878 462604 1878 462604 0 io_out[28]
rlabel metal3 2016 410516 2016 410516 0 io_out[29]
rlabel metal3 581954 99484 581954 99484 0 io_out[2]
rlabel metal3 1832 358428 1832 358428 0 io_out[30]
rlabel metal3 1832 306204 1832 306204 0 io_out[31]
rlabel metal3 1832 254116 1832 254116 0 io_out[32]
rlabel metal2 230874 450286 230874 450286 0 io_out[33]
rlabel metal3 2062 149804 2062 149804 0 io_out[34]
rlabel metal3 475 97580 475 97580 0 io_out[35]
rlabel metal3 1832 58548 1832 58548 0 io_out[36]
rlabel metal3 1924 19380 1924 19380 0 io_out[37]
rlabel metal3 582046 139332 582046 139332 0 io_out[3]
rlabel metal3 582000 179180 582000 179180 0 io_out[4]
rlabel metal3 582092 219028 582092 219028 0 io_out[5]
rlabel metal2 579830 259131 579830 259131 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 365381 580198 365381 0 io_out[8]
rlabel metal2 580198 418863 580198 418863 0 io_out[9]
rlabel metal2 194665 250036 194665 250036 0 la_data_in[0]
rlabel metal2 197478 132236 197478 132236 0 la_data_out[0]
rlabel metal2 481758 2030 481758 2030 0 la_data_out[100]
rlabel metal2 485254 2047 485254 2047 0 la_data_out[101]
rlabel metal2 488842 2812 488842 2812 0 la_data_out[102]
rlabel metal2 339565 250036 339565 250036 0 la_data_out[103]
rlabel metal2 495926 2778 495926 2778 0 la_data_out[104]
rlabel metal2 342325 250036 342325 250036 0 la_data_out[105]
rlabel metal2 503010 2744 503010 2744 0 la_data_out[106]
rlabel metal2 506506 2710 506506 2710 0 la_data_out[107]
rlabel metal2 346465 250036 346465 250036 0 la_data_out[108]
rlabel metal2 347898 249009 347898 249009 0 la_data_out[109]
rlabel metal2 211225 250036 211225 250036 0 la_data_out[10]
rlabel metal2 349225 250036 349225 250036 0 la_data_out[110]
rlabel metal2 350605 250036 350605 250036 0 la_data_out[111]
rlabel metal2 351985 250036 351985 250036 0 la_data_out[112]
rlabel metal2 353418 248669 353418 248669 0 la_data_out[113]
rlabel metal1 357006 98668 357006 98668 0 la_data_out[114]
rlabel metal3 356707 247180 356707 247180 0 la_data_out[115]
rlabel metal2 538430 3254 538430 3254 0 la_data_out[116]
rlabel metal2 542018 3951 542018 3951 0 la_data_out[117]
rlabel metal2 545514 4648 545514 4648 0 la_data_out[118]
rlabel metal2 361645 250036 361645 250036 0 la_data_out[119]
rlabel metal2 212658 248176 212658 248176 0 la_data_out[11]
rlabel metal2 363025 250036 363025 250036 0 la_data_out[120]
rlabel metal2 364405 250036 364405 250036 0 la_data_out[121]
rlabel metal2 365785 250036 365785 250036 0 la_data_out[122]
rlabel metal2 367165 250036 367165 250036 0 la_data_out[123]
rlabel metal2 368598 246782 368598 246782 0 la_data_out[124]
rlabel metal2 369925 250036 369925 250036 0 la_data_out[125]
rlabel metal2 371358 246102 371358 246102 0 la_data_out[126]
rlabel metal2 372685 250036 372685 250036 0 la_data_out[127]
rlabel metal2 213985 250036 213985 250036 0 la_data_out[12]
rlabel metal2 172953 340 172953 340 0 la_data_out[13]
rlabel metal2 176686 121268 176686 121268 0 la_data_out[14]
rlabel metal2 218125 250036 218125 250036 0 la_data_out[15]
rlabel metal1 201526 102782 201526 102782 0 la_data_out[16]
rlabel metal2 187121 340 187121 340 0 la_data_out[17]
rlabel metal2 190854 1962 190854 1962 0 la_data_out[18]
rlabel metal2 194442 1996 194442 1996 0 la_data_out[19]
rlabel metal2 198805 250036 198805 250036 0 la_data_out[1]
rlabel metal2 197938 3627 197938 3627 0 la_data_out[20]
rlabel metal2 201526 3627 201526 3627 0 la_data_out[21]
rlabel metal2 205114 1894 205114 1894 0 la_data_out[22]
rlabel metal2 229218 248737 229218 248737 0 la_data_out[23]
rlabel metal2 211961 340 211961 340 0 la_data_out[24]
rlabel metal2 215503 340 215503 340 0 la_data_out[25]
rlabel metal1 232254 247078 232254 247078 0 la_data_out[26]
rlabel metal2 217442 132974 217442 132974 0 la_data_out[27]
rlabel metal2 236118 249196 236118 249196 0 la_data_out[28]
rlabel metal2 229862 1826 229862 1826 0 la_data_out[29]
rlabel metal2 134182 1962 134182 1962 0 la_data_out[2]
rlabel metal2 233450 1860 233450 1860 0 la_data_out[30]
rlabel metal2 237038 2234 237038 2234 0 la_data_out[31]
rlabel metal2 240534 2200 240534 2200 0 la_data_out[32]
rlabel metal2 244122 2166 244122 2166 0 la_data_out[33]
rlabel metal2 247618 2132 247618 2132 0 la_data_out[34]
rlabel metal2 251206 2098 251206 2098 0 la_data_out[35]
rlabel metal2 254702 2064 254702 2064 0 la_data_out[36]
rlabel metal2 248538 248924 248538 248924 0 la_data_out[37]
rlabel metal2 249918 248856 249918 248856 0 la_data_out[38]
rlabel metal2 251245 250036 251245 250036 0 la_data_out[39]
rlabel metal2 137678 1996 137678 1996 0 la_data_out[3]
rlabel metal2 252625 250036 252625 250036 0 la_data_out[40]
rlabel metal2 272458 1894 272458 1894 0 la_data_out[41]
rlabel metal2 255385 250036 255385 250036 0 la_data_out[42]
rlabel metal2 256818 248941 256818 248941 0 la_data_out[43]
rlabel metal2 283130 1979 283130 1979 0 la_data_out[44]
rlabel metal2 259525 250036 259525 250036 0 la_data_out[45]
rlabel metal2 290214 1843 290214 1843 0 la_data_out[46]
rlabel metal2 293710 3356 293710 3356 0 la_data_out[47]
rlabel metal2 263665 250036 263665 250036 0 la_data_out[48]
rlabel metal2 300794 3322 300794 3322 0 la_data_out[49]
rlabel metal2 141266 1894 141266 1894 0 la_data_out[4]
rlabel metal2 266425 250036 266425 250036 0 la_data_out[50]
rlabel metal2 307970 1894 307970 1894 0 la_data_out[51]
rlabel metal2 269185 250036 269185 250036 0 la_data_out[52]
rlabel metal2 270565 250036 270565 250036 0 la_data_out[53]
rlabel metal2 271998 248856 271998 248856 0 la_data_out[54]
rlabel metal2 273325 250036 273325 250036 0 la_data_out[55]
rlabel metal2 274705 250036 274705 250036 0 la_data_out[56]
rlabel metal2 329222 2098 329222 2098 0 la_data_out[57]
rlabel metal2 332718 2132 332718 2132 0 la_data_out[58]
rlabel metal2 278845 250036 278845 250036 0 la_data_out[59]
rlabel metal2 179262 125834 179262 125834 0 la_data_out[5]
rlabel metal2 280225 250036 280225 250036 0 la_data_out[60]
rlabel metal2 281605 250036 281605 250036 0 la_data_out[61]
rlabel metal2 346978 1860 346978 1860 0 la_data_out[62]
rlabel metal2 350474 1826 350474 1826 0 la_data_out[63]
rlabel metal2 354062 1792 354062 1792 0 la_data_out[64]
rlabel metal2 287125 250036 287125 250036 0 la_data_out[65]
rlabel metal2 288505 250036 288505 250036 0 la_data_out[66]
rlabel metal1 290904 247078 290904 247078 0 la_data_out[67]
rlabel metal2 367993 340 367993 340 0 la_data_out[68]
rlabel metal2 371489 340 371489 340 0 la_data_out[69]
rlabel metal2 148350 1928 148350 1928 0 la_data_out[6]
rlabel metal1 295044 247078 295044 247078 0 la_data_out[70]
rlabel metal2 295405 250036 295405 250036 0 la_data_out[71]
rlabel metal1 340538 232526 340538 232526 0 la_data_out[72]
rlabel metal2 385526 16560 385526 16560 0 la_data_out[73]
rlabel metal2 389344 16560 389344 16560 0 la_data_out[74]
rlabel metal2 392833 340 392833 340 0 la_data_out[75]
rlabel metal2 302305 250036 302305 250036 0 la_data_out[76]
rlabel metal2 303685 250036 303685 250036 0 la_data_out[77]
rlabel metal2 403328 16560 403328 16560 0 la_data_out[78]
rlabel metal2 306498 248992 306498 248992 0 la_data_out[79]
rlabel metal2 151846 2064 151846 2064 0 la_data_out[7]
rlabel metal2 307878 248958 307878 248958 0 la_data_out[80]
rlabel metal2 309258 248924 309258 248924 0 la_data_out[81]
rlabel metal2 310585 250036 310585 250036 0 la_data_out[82]
rlabel metal2 312018 249094 312018 249094 0 la_data_out[83]
rlabel metal2 424994 1758 424994 1758 0 la_data_out[84]
rlabel metal2 314778 249162 314778 249162 0 la_data_out[85]
rlabel metal2 316158 249128 316158 249128 0 la_data_out[86]
rlabel metal2 317485 250036 317485 250036 0 la_data_out[87]
rlabel metal2 318865 250036 318865 250036 0 la_data_out[88]
rlabel metal2 442658 7402 442658 7402 0 la_data_out[89]
rlabel metal2 155434 2098 155434 2098 0 la_data_out[8]
rlabel metal2 446246 1860 446246 1860 0 la_data_out[90]
rlabel metal2 449834 2234 449834 2234 0 la_data_out[91]
rlabel metal2 324385 250036 324385 250036 0 la_data_out[92]
rlabel metal2 325818 247462 325818 247462 0 la_data_out[93]
rlabel metal2 327145 250036 327145 250036 0 la_data_out[94]
rlabel metal2 328525 250036 328525 250036 0 la_data_out[95]
rlabel metal2 329905 250036 329905 250036 0 la_data_out[96]
rlabel metal2 331338 248788 331338 248788 0 la_data_out[97]
rlabel metal2 332718 246816 332718 246816 0 la_data_out[98]
rlabel metal2 334045 250036 334045 250036 0 la_data_out[99]
rlabel metal2 209845 250036 209845 250036 0 la_data_out[9]
rlabel metal1 195684 247078 195684 247078 0 la_oenb[0]
rlabel metal3 156588 99216 156588 99216 0 low
rlabel metal2 334926 498790 334926 498790 0 reset
rlabel metal2 370070 680891 370070 680891 0 start
rlabel metal2 271998 681231 271998 681231 0 uP_data_mem_addr\[0\]
rlabel metal2 274390 681163 274390 681163 0 uP_data_mem_addr\[1\]
rlabel metal2 276782 681214 276782 681214 0 uP_data_mem_addr\[2\]
rlabel metal2 195086 591396 195086 591396 0 uP_data_mem_addr\[3\]
rlabel metal2 281566 681146 281566 681146 0 uP_data_mem_addr\[4\]
rlabel metal2 283958 681027 283958 681027 0 uP_data_mem_addr\[5\]
rlabel metal2 286350 681095 286350 681095 0 uP_data_mem_addr\[6\]
rlabel metal2 288742 680959 288742 680959 0 uP_data_mem_addr\[7\]
rlabel metal2 367678 681163 367678 681163 0 uP_dataw_en
rlabel metal1 218454 496230 218454 496230 0 uP_instr\[0\]
rlabel via1 250102 679405 250102 679405 0 uP_instr\[10\]
rlabel metal2 255017 449956 255017 449956 0 uP_instr\[11\]
rlabel metal2 256489 449956 256489 449956 0 uP_instr\[12\]
rlabel metal4 264500 678980 264500 678980 0 uP_instr\[13\]
rlabel metal2 267214 680364 267214 680364 0 uP_instr\[14\]
rlabel metal4 269284 678912 269284 678912 0 uP_instr\[15\]
rlabel metal1 219006 460666 219006 460666 0 uP_instr\[1\]
rlabel metal1 219328 462910 219328 462910 0 uP_instr\[2\]
rlabel metal2 216982 680908 216982 680908 0 uP_instr\[3\]
rlabel metal2 221766 681282 221766 681282 0 uP_instr\[4\]
rlabel metal2 226550 681112 226550 681112 0 uP_instr\[5\]
rlabel metal2 231334 681078 231334 681078 0 uP_instr\[6\]
rlabel metal2 236118 681044 236118 681044 0 uP_instr\[7\]
rlabel metal2 195822 572662 195822 572662 0 uP_instr\[8\]
rlabel metal2 251390 463445 251390 463445 0 uP_instr\[9\]
rlabel metal2 236210 461881 236210 461881 0 uP_instr_mem_addr\[0\]
rlabel metal2 254111 449956 254111 449956 0 uP_instr_mem_addr\[10\]
rlabel metal2 257646 680432 257646 680432 0 uP_instr_mem_addr\[11\]
rlabel metal2 256857 449956 256857 449956 0 uP_instr_mem_addr\[12\]
rlabel metal1 218408 465562 218408 465562 0 uP_instr_mem_addr\[1\]
rlabel metal1 220892 465630 220892 465630 0 uP_instr_mem_addr\[2\]
rlabel metal2 219374 680874 219374 680874 0 uP_instr_mem_addr\[3\]
rlabel metal2 195730 572900 195730 572900 0 uP_instr_mem_addr\[4\]
rlabel metal2 195638 572798 195638 572798 0 uP_instr_mem_addr\[5\]
rlabel metal2 233726 681010 233726 681010 0 uP_instr_mem_addr\[6\]
rlabel metal2 238510 681299 238510 681299 0 uP_instr_mem_addr\[7\]
rlabel metal1 223652 468622 223652 468622 0 uP_instr_mem_addr\[8\]
rlabel metal1 227010 468690 227010 468690 0 uP_instr_mem_addr\[9\]
rlabel metal2 215694 500412 215694 500412 0 uP_read_data\[0\]
rlabel metal2 315054 680194 315054 680194 0 uP_read_data\[10\]
rlabel metal2 255898 450932 255898 450932 0 uP_read_data\[11\]
rlabel metal2 257370 450966 257370 450966 0 uP_read_data\[12\]
rlabel metal2 258375 449956 258375 449956 0 uP_read_data\[13\]
rlabel metal1 324898 679218 324898 679218 0 uP_read_data\[14\]
rlabel metal2 327014 681299 327014 681299 0 uP_read_data\[15\]
rlabel metal2 195270 588693 195270 588693 0 uP_read_data\[1\]
rlabel metal2 195362 588387 195362 588387 0 uP_read_data\[2\]
rlabel metal3 296700 679184 296700 679184 0 uP_read_data\[3\]
rlabel metal1 220708 497658 220708 497658 0 uP_read_data\[4\]
rlabel metal2 303094 680330 303094 680330 0 uP_read_data\[5\]
rlabel metal3 199916 576980 199916 576980 0 uP_read_data\[6\]
rlabel metal2 307878 680296 307878 680296 0 uP_read_data\[7\]
rlabel metal2 310270 680262 310270 680262 0 uP_read_data\[8\]
rlabel metal2 312662 680228 312662 680228 0 uP_read_data\[9\]
rlabel metal2 329406 680160 329406 680160 0 uP_write_data\[0\]
rlabel metal2 254649 449956 254649 449956 0 uP_write_data\[10\]
rlabel metal2 256121 449956 256121 449956 0 uP_write_data\[11\]
rlabel metal2 257593 449956 257593 449956 0 uP_write_data\[12\]
rlabel metal2 258697 449956 258697 449956 0 uP_write_data\[13\]
rlabel metal2 259801 449956 259801 449956 0 uP_write_data\[14\]
rlabel metal2 365286 680942 365286 680942 0 uP_write_data\[15\]
rlabel metal2 331798 680143 331798 680143 0 uP_write_data\[1\]
rlabel metal2 334190 681282 334190 681282 0 uP_write_data\[2\]
rlabel metal2 336582 681248 336582 681248 0 uP_write_data\[3\]
rlabel metal4 372692 588472 372692 588472 0 uP_write_data\[4\]
rlabel metal4 373796 588472 373796 588472 0 uP_write_data\[5\]
rlabel metal2 343758 681010 343758 681010 0 uP_write_data\[6\]
rlabel metal2 346150 680976 346150 680976 0 uP_write_data\[7\]
rlabel metal2 348542 681044 348542 681044 0 uP_write_data\[8\]
rlabel metal2 350934 681078 350934 681078 0 uP_write_data\[9\]
rlabel metal2 581026 1724 581026 1724 0 user_irq[0]
rlabel metal2 582222 1894 582222 1894 0 user_irq[1]
rlabel metal2 582912 16560 582912 16560 0 user_irq[2]
rlabel metal2 361 340 361 340 0 wb_clk_i
rlabel metal2 1557 340 1557 340 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
